`define CYCLE_TIME 20.0
`define NUMBER_OF_PAT 100
module PATTERN(
        // Input signals
        clk,
        rst_n,
        i_valid,
        w_valid,
        i_data,
        w_data,
        // Output signals
        w_ready,
        o_valid,
        o_data
);
//================================================================
// I/O PORTS
//================================================================
output logic clk, rst_n, i_valid, w_valid;
output logic [7:0] i_data, w_data;

input w_ready, o_valid;
input [31:0] o_data;
//================================================================
// wire & registers
//================================================================
logic  [7:0] i_mtx   [0:7][0:15];
logic  [7:0] i_t_mtx [0:15][0:7];
logic [23:0] a_mtx   [0:7][0:7];
logic  [7:0] w_mtx   [0:7];
logic [31:0] o_mtx   [0:7];
logic [31:0] sum     [0:7];
logic [31:0] avg     [0:7];
//================================================================
// PARAMETERS & VARIABLES
//================================================================
integer i, j, k;
integer PATNUM, patcount;
integer pat_delay, input_gap;
integer lat, lat_check, latency;
integer w_ready_cnt, o_valid_cnt, ready_cnt;
real	CYCLE = `CYCLE_TIME;
always	#(CYCLE/2.0) clk = ~clk;
//================================================================
// SPEC 3 : Check i_valid and w_ready overlap or not
//================================================================
always @ (*) begin 
	if (w_ready === 1 && i_valid === 1) begin 
		fail ;
		$display ("-------------------------------------------------------------------------------------------------------------------------------------");
		$display ("                                                       FAIL!                                                                         ");
		$display ("                                               SPEC 3 is violated                                                                    ");
		$display ("                                         i_valid and w_ready cannot be overlapped                                                    ");
		$display ("-------------------------------------------------------------------------------------------------------------------------------------");
		$finish ;
	end
end
//================================================================
// SPEC 5 : Check w_valid and o_valid overlap or not
//================================================================
always @ (*) begin 
	if (o_valid === 1 && w_valid === 1) begin 
		fail ;
		$display ("-------------------------------------------------------------------------------------------------------------------------------------");
		$display ("                                                       FAIL!                                                                         ");
		$display ("                                               SPEC 5 is violated                                                                    ");
		$display ("                                         w_valid and o_valid cannot be overlapped                                                    ");
		$display ("-------------------------------------------------------------------------------------------------------------------------------------");
		$finish ;
	end
end
//================================================================
// SPEC 7 : Check all output should be reset when o_valid is low
//================================================================
always @ (negedge clk) begin
	if (o_valid === 0 && o_data !== 0) begin
		fail ;
		$display ("-------------------------------------------------------------------------------------------------------------------------------------");
		$display ("                                                       FAIL!                                                                         ");
		$display ("                                               SPEC 7 is violated                                                                    ");
		$display ("                                        All outputs should be zero when o_valid is low                                               ");
		$display ("-------------------------------------------------------------------------------------------------------------------------------------");
		$finish ;	
	end
end
//================================================================
// w_ready could be pulled high once for each pat_number
//================================================================
always @ (negedge clk) begin
	if (w_ready) begin
		ready_cnt = ready_cnt + 1;
	end
end
//================================================================
// initial
//================================================================
initial begin
	latency = 0;
	ready_cnt = -1;
	rst_n = 1'b1;
	i_valid = 0;
	w_valid = 0;
	i_data = 'bx;
	w_data = 'bx;

	force clk = 0;
	RESET_TASK;
	PATNUM = `NUMBER_OF_PAT;
	for(patcount = 0; patcount < PATNUM; patcount = patcount + 1) begin
		pat_delay = $urandom_range(5,10) ;
		repeat(pat_delay) @(negedge clk) ;
		INPUT_TASK;
		WAIT_W_READY;
		CHECK_W_READY;
		WEIGHT_TASK;
		WAIT_O_VALID;
		CHECK_ANS;
		case(patcount % 5)
		0 : $display("\033[31m PASS PATTERN NO.%3d", patcount);
		1 : $display("\033[32m PASS PATTERN NO.%3d", patcount);
		2 : $display("\033[33m PASS PATTERN NO.%3d", patcount);
		3 : $display("\033[34m PASS PATTERN NO.%3d", patcount);
		4 : $display("\033[35m PASS PATTERN NO.%3d", patcount);
		endcase
		$display(" The execution latency of PATTERN NO.%3d is %3d", patcount, lat);
		if(patcount !== ready_cnt)begin
			fail ;
			$display ("-------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                       FAIL!                                                                         ");
			$display ("                                   w_ready could be pulled high once for each pat_number                                             ");
			$display ("-------------------------------------------------------------------------------------------------------------------------------------");
			$finish ;				
		end
	end
	YOU_PASS_task;

	$finish;
end

//================================================================
// task
//================================================================
task RESET_TASK; begin
    #(CYCLE); rst_n = 0;
    #(CYCLE);
    if(w_ready !== 0 || o_valid !== 0 || o_data !== 0) begin
        fail;
	    $display ("-------------------------------------------------------------------------------------------------------------------------------------");
		$display ("                                                              FAIL!                                                                  ");
		$display ("                                                       SPEC 2 is violated                                                            ");
		$display ("                                              All outputs should be 0 after reset                                                    ");
		$display ("-------------------------------------------------------------------------------------------------------------------------------------");
		$finish ;
    end
	rst_n = 1 ;
    #(20); release clk;	
end endtask

task INPUT_TASK; begin
    i_valid = 1;
	lat = 0;
	for (i = 0 ; i < 8 ; i = i + 1) begin
		for (j = 0 ; j < 16 ; j = j + 1) begin
			lat = lat + 1;
			i_mtx[i][j] = $urandom_range(0,255);
			i_t_mtx[j][i] = i_mtx[i][j];
			i_data = i_mtx[i][j];
			@(negedge clk);
		end
	end
	i_valid = 0;
	i_data = 'bx;
	lat_check = -1;
end endtask

task WAIT_W_READY; begin
	while (w_ready !== 1) begin
		lat = lat + 1;
		lat_check = lat_check + 1;
        if(lat_check == 10000) begin
			fail ;
			$display ("-------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                              FAIL!                                                                  ");
			$display ("                                                        SPEC 4 is violated                                                           ");
			$display ("                                              The w_ready signal hasn't been received                                                ");
			$display ("                                                         Pattern No. %3d                                                             ", patcount);
			$display ("                                             The execution latency are over 1000 cycles                                              ");
			$display ("-------------------------------------------------------------------------------------------------------------------------------------");
			repeat(2) @(negedge clk) ;
			$finish ;
        end
	@(negedge clk) ;
	end
	// MM 1
	for (i = 0 ; i < 8 ; i = i + 1) begin
		for (j = 0 ; j < 8 ; j = j + 1) begin
			a_mtx[i][j] = 0;
			for (k = 0 ; k < 16 ; k = k + 1) begin
				a_mtx[i][j] = a_mtx[i][j] + i_mtx[i][k] * i_t_mtx[k][j];
			end
		end
	end
	// RAT
	for (i = 0 ; i < 8 ; i = i + 1) begin
		sum[i] = 0;
		avg[i] = 0;
		for (j = 0 ; j < 8 ; j = j + 1) begin
			sum[i] = sum[i] + a_mtx[i][j];
		end
		avg[i] = sum[i] / 8;
	end
	for (i = 0 ; i < 8 ; i = i + 1) begin
		for (j = 0 ; j < 8 ; j = j + 1) begin
			if (a_mtx[i][j] < avg[i]) begin
				a_mtx[i][j] = 0;
			end
			else begin
				a_mtx[i][j] = a_mtx[i][j];
			end
		end
	end
end endtask

task CHECK_W_READY; begin
	w_ready_cnt = 0;
    while(w_ready === 1) begin
		lat = lat + 1;
		lat_check = lat_check + 1;
        if(w_ready_cnt == 1) begin
            fail;
            $display ("-------------------------------------------------------------------------------------------------------------------------------------");
            $display ("                                                                FAIL !                                                               ");
			$display ("                                                         Pattern No. %3d                                                             ", patcount);
            $display ("                                               w_ready should be pulled high for only 1 cycle!                                       ");
            $display ("-------------------------------------------------------------------------------------------------------------------------------------");
			#(100);
			$finish;
        end
		w_ready_cnt = w_ready_cnt + 1;		
        @(negedge clk);
    end
	if(w_ready_cnt !== 1) begin
		fail;
		$display ("-------------------------------------------------------------------------------------------------------------------------------------");
		$display ("                                                                FAIL !                                                               ");
		$display ("                                                         Pattern No. %3d                                                             ", patcount);
		$display ("                                               w_ready should be pulled high for only 1 cycle!                                       ");
		$display ("-------------------------------------------------------------------------------------------------------------------------------------");
		#(100);
		$finish;
	end
	w_ready_cnt = 0;
end endtask

task WEIGHT_TASK; begin
    input_gap = $urandom_range(2,6);
    repeat(input_gap) @(negedge clk);
	lat = lat + input_gap;
	lat_check = lat_check + input_gap;
    w_valid = 1;
    for(i = 0; i < 8; i = i + 1) begin
		lat = lat + 1;
		lat_check = lat_check + 1;
		w_mtx[i] = $urandom_range(0,255);
		w_data = w_mtx[i];
		@(negedge clk);
	end
	w_valid = 0;
	w_data = 'bx;
	// MM2
	for (i = 0 ; i < 8 ; i = i + 1) begin
		o_mtx[i] = 0;
		for (j = 0 ; j < 8 ; j = j + 1) begin
			o_mtx[i] = o_mtx[i] + a_mtx[i][j] * w_mtx[j];
		end
	end
end endtask

task WAIT_O_VALID; begin
    while(o_valid !== 1) begin
        lat = lat + 1;
		lat_check = lat_check + 1;
        if(lat_check == 10000) begin
			fail ;
			$display ("-------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                              FAIL!                                                                  ");
			$display ("                                                        SPEC 4 is violated                                                           ");
			$display ("                                              The o_valid signal hasn't been received                                                ");
			$display ("                                                         Pattern No. %3d                                                             ", patcount);
			$display ("                                             The execution latency are over 1000 cycles                                              ");
			$display ("-------------------------------------------------------------------------------------------------------------------------------------");
			repeat(2) @(negedge clk) ;
			$finish ;
        end
        @(negedge clk);
    end
end endtask

task CHECK_ANS ; begin
	o_valid_cnt = 0;
	while(o_valid === 1) begin
		lat = lat + 1;
		lat_check = lat_check + 1;
		if(o_valid_cnt === 8)begin
			fail;
			$display ("-------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                              FAIL!                                                                  ");
			$display ("                                                        SPEC 6 is violated                                                           ");
			$display ("                                                         Pattern No. %3d                                                             ", patcount);
			$display ("                                                Output should be output only for 8 cycles                                             ");
			$display ("-------------------------------------------------------------------------------------------------------------------------------------");
			#(100);
			$finish ;		
		end
		if (o_data !== o_mtx[o_valid_cnt]) begin
			fail;
			$display ("-------------------------------------------------------------------------------------------------------------------------------------");
			$display ("                                                               FAIL!                                                                 ");
			$display ("                                                         Pattern No. %3d                                                             ", patcount);
			$display ("                                         ERROR occurs at the %3d th element of the output vector                                     ", o_valid_cnt);
			$display ("                                                         YOUR answer : %d                                                            ",o_data);
			$display ("                                                       GOLDEN answer : %d                                                            ",o_mtx[o_valid_cnt]);
			$display ("-------------------------------------------------------------------------------------------------------------------------------------");
			#(100);
			$finish;			
		end
		o_valid_cnt = o_valid_cnt + 1;
		@(negedge clk);
	end
	latency = latency + lat;
	if(o_valid_cnt !== 8)begin
		fail;
		$display ("-------------------------------------------------------------------------------------------------------------------------------------");
		$display ("                                                              FAIL!                                                                  ");
		$display ("                                                        SPEC 6 is violated                                                           ");
		$display ("                                                         Pattern No. %3d                                                             ", patcount);
		$display ("                                                Output should be output only for 8 cycles                                             ");
		$display ("-------------------------------------------------------------------------------------------------------------------------------------");
		#(100);
		$finish ;		
	end
	o_valid_cnt = 0;
end endtask

task YOU_PASS_task;begin
$display("\033[37m                                                                                                                                          ");        
$display("\033[37m                                                                                \033[32m      :BBQvi.                                              ");        
$display("\033[37m                                                              .i7ssrvs7         \033[32m     BBBBBBBBQi                                           ");        
$display("\033[37m                        .:r7rrrr:::.        .::::::...   .i7vr:.      .B:       \033[32m    :BBBP :7BBBB.                                         ");        
$display("\033[37m                      .Kv.........:rrvYr7v7rr:.....:rrirJr.   .rgBBBBg  Bi      \033[32m    BBBB     BBBB                                         ");        
$display("\033[37m                     7Q  :rubEPUri:.       ..:irrii:..    :bBBBBBBBBBBB  B      \033[32m   iBBBv     BBBB       vBr                               ");        
$display("\033[37m                    7B  BBBBBBBBBBBBBBB::BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB :R     \033[32m   BBBBBKrirBBBB.     :BBBBBB:                            ");        
$display("\033[37m                   Jd .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: Bi    \033[32m  rBBBBBBBBBBBR.    .BBBM:BBB                             ");        
$display("\033[37m                  uZ .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB .B    \033[32m  BBBB   .::.      EBBBi :BBU                             ");        
$display("\033[37m                 7B .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  B    \033[32m MBBBr           vBBBu   BBB.                             ");        
$display("\033[37m                .B  BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: JJ   \033[32m i7PB          iBBBBB.  iBBB                              ");        
$display("\033[37m                B. BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  Lu             \033[32m  vBBBBPBBBBPBBB7       .7QBB5i                ");        
$display("\033[37m               Y1 KBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBi XBBBBBBBi :B            \033[32m :RBBB.  .rBBBBB.      rBBBBBBBB7              ");        
$display("\033[37m              :B .BBBBBBBBBBBBBsRBBBBBBBBBBBrQBBBBB. UBBBRrBBBBBBr 1BBBBBBBBB  B.          \033[32m    .       BBBB       BBBB  :BBBB             ");        
$display("\033[37m              Bi BBBBBBBBBBBBBi :BBBBBBBBBBE .BBK.  .  .   QBBBBBBBBBBBBBBBBBB  Bi         \033[32m           rBBBr       BBBB    BBBU            ");        
$display("\033[37m             .B .BBBBBBBBBBBBBBQBBBBBBBBBBBB       \033[38;2;242;172;172mBBv \033[37m.LBBBBBBBBBBBBBBBBBBBBBB. B7.:ii:   \033[32m           vBBB        .BBBB   :7i.            ");        
$display("\033[37m            .B  PBBBBBBBBBBBBBBBBBBBBBBBBBBBBbYQB. \033[38;2;242;172;172mBB: \033[37mBBBBBBBBBBBBBBBBBBBBBBBBB  Jr:::rK7 \033[32m             .7  BBB7   iBBBg                  ");        
$display("\033[37m           7M  PBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  \033[38;2;242;172;172mBB. \033[37mBBBBBBBBBBBBBBBBBBBBBBB..i   .   v1                  \033[32mdBBB.   5BBBr                 ");        
$display("\033[37m          sZ .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  \033[38;2;242;172;172mBB. \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBB iD2BBQL.                 \033[32m ZBBBr  EBBBv     YBBBBQi     ");        
$display("\033[37m  .7YYUSIX5 .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  \033[38;2;242;172;172mBB. \033[37mBBBBBBBBBBBBBBBBBBBBBBBBY.:.      :B                 \033[32m  iBBBBBBBBD     BBBBBBBBB.   ");        
$display("\033[37m LB.        ..BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB. \033[38;2;242;172;172mBB: \033[37mBBBBBBBBBBBBBBBBBBBBBBBBMBBB. BP17si                 \033[32m    :LBBBr      vBBBi  5BBB   ");        
$display("\033[37m  KvJPBBB :BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: \033[38;2;242;172;172mZB: \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBsiJr .i7ssr:                \033[32m          ...   :BBB:   BBBu  ");        
$display("\033[37m i7ii:.   ::BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBj \033[38;2;242;172;172muBi \033[37mQBBBBBBBBBBBBBBBBBBBBBBBBi.ir      iB                \033[32m         .BBBi   BBBB   iMBu  ");        
$display("\033[37mDB    .  vBdBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBg \033[38;2;242;172;172m7Bi \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBBBB rBrXPv.                \033[32m          BBBX   :BBBr        ");        
$display("\033[37m :vQBBB. BQBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBQ \033[38;2;242;172;172miB: \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBBBB .L:ii::irrrrrrrr7jIr   \033[32m          .BBBv  :BBBQ        ");        
$display("\033[37m :7:.   .. 5BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  \033[38;2;242;172;172mBr \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBBB:            ..... ..YB. \033[32m           .BBBBBBBBB:        ");        
$display("\033[37mBU  .:. BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  \033[38;2;242;172;172mB7 \033[37mgBBBBBBBBBBBBBBBBBBBBBBBBBB. gBBBBBBBBBBBBBBBBBB. BL \033[32m             rBBBBB1.         ");        
$display("\033[37m rY7iB: BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: \033[38;2;242;172;172mB7 \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBB. QBBBBBBBBBBBBBBBBBi  v5                                ");        
$display("\033[37m     us EBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB \033[38;2;242;172;172mIr \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBgu7i.:BBBBBBBr Bu                                 ");        
$display("\033[37m      B  7BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB.\033[38;2;242;172;172m:i \033[37mBBBBBBBBBBBBBBBBBBBBBBBBBBBv:.  .. :::  .rr    rB                                  ");        
$display("\033[37m      us  .BBBBBBBBBBBBBQLXBBBBBBBBBBBBBBBBBBBBBBBBq  .BBBBBBBBBBBBBBBBBBBBBBBBBv  :iJ7vri:::1Jr..isJYr                                   ");        
$display("\033[37m      B  BBBBBBB  MBBBM      qBBBBBBBBBBBBBBBBBBBBBB: BBBBBBBBBBBBBBBBBBBBBBBBBB  B:           iir:                                       ");        
$display("\033[37m     iB iBBBBBBBL       BBBP. :BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  B.                                                       ");        
$display("\033[37m     P: BBBBBBBBBBB5v7gBBBBBB  BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: Br                                                        ");        
$display("\033[37m     B  BBBs 7BBBBBBBBBBBBBB7 :BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB .B                                                         ");        
$display("\033[37m    .B :BBBB.  EBBBBBQBBBBBJ .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB. B.                                                         ");        
$display("\033[37m    ij qBBBBBg          ..  .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB .B                                                          ");        
$display("\033[37m    UY QBBBBBBBBSUSPDQL...iBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBK EL                                                          ");        
$display("\033[37m    B7 BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB: B:                                                          ");        
$display("\033[37m    B  BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBYrBB vBBBBBBBBBBBBBBBBBBBBBBBB. Ls                                                          ");        
$display("\033[37m    B  BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBi_  /UBBBBBBBBBBBBBBBBBBBBBBBBB. :B:                                                        ");        
$display("\033[37m   rM .BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB  ..IBBBBBBBBBBBBBBBBQBBBBBBBBBB  B                                                        ");        
$display("\033[37m   B  BBBBBBBBBdZBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBPBBBBBBBBBBBBEji:..     sBBBBBBBr Br                                                       ");        
$display("\033[37m  7B 7BBBBBBBr     .:vXQBBBBBBBBBBBBBBBBBBBBBBBBBQqui::..  ...i:i7777vi  BBBBBBr Bi                                                       ");        
$display("\033[37m  Ki BBBBBBB  rY7vr:i....  .............:.....  ...:rii7vrr7r:..      7B  BBBBB  Bi                                                       ");        
$display("\033[37m  B. BBBBBB  B:    .::ir77rrYLvvriiiiiiirvvY7rr77ri:..                 bU  iQBB:..rI                                                      ");        
$display("\033[37m.S: 7BBBBP  B.                                                          vI7.  .:.  B.                                                     ");        
$display("\033[37mB: ir:.   :B.                                                    ");
$display("\033[35mDofuramingo is the cutest kitty                                                                                                                            \033[m");
$display ("----------------------------------------------------------------------------------------------------------------------");
$display ("                                                  Congratulations!                                                                        ");
$display ("                                           You have passed all patterns!                                                                  ");
$display ("                                           Average Latency : %3f ns                                                                   ", (latency / patcount)*CYCLE);
$display ("                                             cycle time    : %3f ns                                                                     ",CYCLE);
$display ("----------------------------------------------------------------------------------------------------------------------");

$finish;
end endtask

task fail; begin
$display("\033[38;2;252;238;238m                                                                                                                                           ");      
$display("\033[38;2;252;238;238m                                                                                                :L777777v7.                                ");
$display("\033[31m  i:..::::::i.      :::::         ::::    .:::.       \033[38;2;252;238;238m                                       .vYr::::::::i7Lvi                             ");
$display("\033[31m  BBBBBBBBBBBi     iBBBBBL       .BBBB    7BBB7       \033[38;2;252;238;238m                                      JL..\033[38;2;252;172;172m:r777v777i::\033[38;2;252;238;238m.ijL                           ");
$display("\033[31m  BBBB.::::ir.     BBB:BBB.      .BBBv    iBBB:       \033[38;2;252;238;238m                                    :K: \033[38;2;252;172;172miv777rrrrr777v7:.\033[38;2;252;238;238m:J7                         ");
$display("\033[31m  BBBQ            :BBY iBB7       BBB7    :BBB:       \033[38;2;252;238;238m                                   :d \033[38;2;252;172;172m.L7rrrrrrrrrrrrr77v: \033[38;2;252;238;238miI.                       ");
$display("\033[31m  BBBB            BBB. .BBB.      BBB7    :BBB:       \033[38;2;252;238;238m                                  .B \033[38;2;252;172;172m.L7rrrrrrrrrrrrrrrrr7v..\033[38;2;252;238;238mBr                      ");
$display("\033[31m  BBBB:r7vvj:    :BBB   gBBs      BBB7    :BBB:       \033[38;2;252;238;238m                                  S:\033[38;2;252;172;172m v7rrrrrrrrrrrrrrrrrrr7v. \033[38;2;252;238;238mB:                     ");
$display("\033[31m  BBBBBBBBBB7    BBB:   .BBB.     BBB7    :BBB:       \033[38;2;252;238;238m                                 .D \033[38;2;252;172;172mi7rrrrrrr777rrrrrrrrrrr7v. \033[38;2;252;238;238mB.                    ");
$display("\033[31m  BBBB    ..    iBBBBBBBBBBBP     BBB7    :BBB:       \033[38;2;252;238;238m                                 rv\033[38;2;252;172;172m v7rrrrrr7rirv7rrrrrrrrrr7v \033[38;2;252;238;238m:I                    ");
$display("\033[31m  BBBB          BBBBi7vviQBBB.    BBB7    :BBB.       \033[38;2;252;238;238m                                 2i\033[38;2;252;172;172m.v7rrrrrr7i  :v7rrrrrrrrrrvi \033[38;2;252;238;238mB:                   ");
$display("\033[31m  BBBB         rBBB.      BBBQ   .BBBv    iBBB2ir777L7\033[38;2;252;238;238m                                 2i.\033[38;2;252;172;172mv7rrrrrr7v \033[38;2;252;238;238m:..\033[38;2;252;172;172mv7rrrrrrrrr77 \033[38;2;252;238;238mrX                   ");
$display("\033[31m .BBBB        :BBBB       BBBB7  .BBBB    7BBBBBBBBBBB\033[38;2;252;238;238m                                 Yv \033[38;2;252;172;172mv7rrrrrrrv.\033[38;2;252;238;238m.B \033[38;2;252;172;172m.vrrrrrrrrrrL.\033[38;2;252;238;238m:5                   ");
$display("\033[31m  . ..        ....         ...:   ....    ..   .......\033[38;2;252;238;238m                                 .q \033[38;2;252;172;172mr7rrrrrrr7i \033[38;2;252;238;238mPv \033[38;2;252;172;172mi7rrrrrrrrrv.\033[38;2;252;238;238m:S                   ");
$display("\033[38;2;252;238;238m                                                                                        Lr \033[38;2;252;172;172m77rrrrrr77 \033[38;2;252;238;238m:B. \033[38;2;252;172;172mv7rrrrrrrrv.\033[38;2;252;238;238m:S                   ");
$display("\033[38;2;252;238;238m                                                                                         B: \033[38;2;252;172;172m7v7rrrrrv. \033[38;2;252;238;238mBY \033[38;2;252;172;172mi7rrrrrrr7v \033[38;2;252;238;238miK                   ");
$display("\033[38;2;252;238;238m                                                                              .::rriii7rir7. \033[38;2;252;172;172m.r77777vi \033[38;2;252;238;238m7B  \033[38;2;252;172;172mvrrrrrrr7r \033[38;2;252;238;238m2r                   ");
$display("\033[38;2;252;238;238m                                                                       .:rr7rri::......    .     \033[38;2;252;172;172m.:i7s \033[38;2;252;238;238m.B. \033[38;2;252;172;172mv7rrrrr7L..\033[38;2;252;238;238mB                    ");
$display("\033[38;2;252;238;238m                                                        .::7L7rriiiirr77rrrrrrrr72BBBBBBBBBBBBvi:..  \033[38;2;252;172;172m.  \033[38;2;252;238;238mBr \033[38;2;252;172;172m77rrrrrvi \033[38;2;252;238;238mKi                    ");
$display("\033[38;2;252;238;238m                                                    :rv7i::...........    .:i7BBBBQbPPPqPPPdEZQBBBBBr:.\033[38;2;252;238;238m ii \033[38;2;252;172;172mvvrrrrvr \033[38;2;252;238;238mvs                     ");
$display("\033[38;2;252;238;238m                    .S77L.                      .rvi:. ..:r7QBBBBBBBBBBBgri.    .:BBBPqqKKqqqqPPPPPEQBBBZi  \033[38;2;252;172;172m:777vi \033[38;2;252;238;238mvI                      ");
$display("\033[38;2;252;238;238m                    B: ..Jv                   isi. .:rBBBBBQZPPPPqqqPPdERBBBBBi.    :BBRKqqqqqqqqqqqqPKDDBB:  \033[38;2;252;172;172m:7. \033[38;2;252;238;238mJr                       ");
$display("\033[38;2;252;238;238m                   vv SB: iu                rL: .iBBBQEPqqPPqqqqqqqqqqqqqPPPPbQBBB:   .EBQKqqqqqqPPPqqKqPPgBB:  .B:                        ");
$display("\033[38;2;252;238;238m                  :R  BgBL..s7            rU: .qBBEKPqqqqqqqqqqqqqqqqqqqqqqqqqPPPEBBB:   EBEPPPEgQBBQEPqqqqKEBB: .s                        ");
$display("\033[38;2;252;238;238m               .U7.  iBZBBBi :ji         5r .MBQqPqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPKgBB:  .BBBBBdJrrSBBQKqqqqKZB7  I:                      ");
$display("\033[38;2;252;238;238m              v2. :rBBBB: .BB:.ru7:    :5. rBQqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPPBB:  :.        .5BKqqqqqqBB. Kr                     ");
$display("\033[38;2;252;238;238m             .B .BBQBB.   .RBBr  :L77ri2  BBqPqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPbBB   \033[38;2;252;172;172m.irrrrri  \033[38;2;252;238;238mQQqqqqqqKRB. 2i                    ");
$display("\033[38;2;252;238;238m              27 :BBU  rBBBdB \033[38;2;252;172;172m iri::::: \033[38;2;252;238;238m.BQKqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqKRBs\033[38;2;252;172;172mirrr7777L: \033[38;2;252;238;238m7BqqqqqqqXZB. BLv772i              ");
$display("\033[38;2;252;238;238m               rY  PK  .:dPMB \033[38;2;252;172;172m.Y77777r.\033[38;2;252;238;238m:BEqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPPBqi\033[38;2;252;172;172mirrrrrv: \033[38;2;252;238;238muBqqqqqqqqqgB  :.:. B:             ");
$display("\033[38;2;252;238;238m                iu 7BBi  rMgB \033[38;2;252;172;172m.vrrrrri\033[38;2;252;238;238mrBEqKqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPQgi\033[38;2;252;172;172mirrrrv. \033[38;2;252;238;238mQQqqqqqqqqqXBb .BBB .s:.           ");
$display("\033[38;2;252;238;238m                i7 BBdBBBPqbB \033[38;2;252;172;172m.vrrrri\033[38;2;252;238;238miDgPPbPqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPQDi\033[38;2;252;172;172mirr77 \033[38;2;252;238;238m:BdqqqqqqqqqqPB. rBB. .:iu7         ");
$display("\033[38;2;252;238;238m                iX.:iBRKPqKXB.\033[38;2;252;172;172m 77rrr\033[38;2;252;238;238mi7QPBBBBPqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPB7i\033[38;2;252;172;172mrr7r \033[38;2;252;238;238m.vBBPPqqqqqqKqBZ  BPBgri: 1B        ");
$display("\033[38;2;252;238;238m                 ivr .BBqqKXBi \033[38;2;252;172;172mr7rri\033[38;2;252;238;238miQgQi   QZKqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPEQi\033[38;2;252;172;172mirr7r.  \033[38;2;252;238;238miBBqPqqqqqqPB:.QPPRBBB LK        ");
$display("\033[38;2;252;238;238m                   :I. iBgqgBZ \033[38;2;252;172;172m:7rr\033[38;2;252;238;238miJQPB.   gRqqqqqqqqPPPPPPPPqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqPQ7\033[38;2;252;172;172mirrr7vr.  \033[38;2;252;238;238mUBqqPPgBBQPBBKqqqKB  B         ");
$display("\033[38;2;252;238;238m                     v7 .BBR: \033[38;2;252;172;172m.r7ri\033[38;2;252;238;238miggqPBrrBBBBBBBBBBBBBBBBBBQEPPqqPPPqqqqqqqqqqqqqqqqqqqqqqqqqPgPi\033[38;2;252;172;172mirrrr7v7  \033[38;2;252;238;238mrBPBBP:.LBbPqqqqqB. u.        ");
$display("\033[38;2;252;238;238m                      .j. . \033[38;2;252;172;172m :77rr\033[38;2;252;238;238miiBPqPbBB::::::.....:::iirrSBBBBBBBQZPPPPPqqqqqqqqqqqqqqqqqqqqEQi\033[38;2;252;172;172mirrrrrr7v \033[38;2;252;238;238m.BB:     :BPqqqqqDB .B        ");
$display("\033[38;2;252;238;238m                       YL \033[38;2;252;172;172m.i77rrrr\033[38;2;252;238;238miLQPqqKQJ. \033[38;2;252;172;172m ............       \033[38;2;252;238;238m..:irBBBBBBZPPPqqqqqqqPPBBEPqqqdRr\033[38;2;252;172;172mirrrrrr7v \033[38;2;252;238;238m.B  .iBB  dQPqqqqPBi Y:       ");
$display("\033[38;2;252;238;238m                     :U:.\033[38;2;252;172;172mrv7rrrrri\033[38;2;252;238;238miPgqqqqKZB.\033[38;2;252;172;172m.v77777777777777ri::..   \033[38;2;252;238;238m  ..:rBBBBQPPqqqqPBUvBEqqqPRr\033[38;2;252;172;172mirrrrrrvi\033[38;2;252;238;238m iB:RBBbB7 :BQqPqKqBR r7       ");
$display("\033[38;2;252;238;238m                    iI.\033[38;2;252;172;172m.v7rrrrrrri\033[38;2;252;238;238midgqqqqqKB:\033[38;2;252;172;172m 77rrrrrrrrrrrrr77777777ri:..   \033[38;2;252;238;238m .:1BBBEPPB:   BbqqPQr\033[38;2;252;172;172mirrrr7vr\033[38;2;252;238;238m .BBBZPqqDB  .JBbqKPBi vi       ");
$display("\033[38;2;252;238;238m                   :B \033[38;2;252;172;172miL7rrrrrrrri\033[38;2;252;238;238mibgqqqqqqBr\033[38;2;252;172;172m r7rrrrrrrrrrrrrrrrrrrrr777777ri:.  \033[38;2;252;238;238m .iBBBBi  .BbqqdRr\033[38;2;252;172;172mirr7v7: \033[38;2;252;238;238m.Bi.dBBPqqgB:  :BPqgB  B        ");
$display("\033[38;2;252;238;238m                   .K.i\033[38;2;252;172;172mv7rrrrrrrri\033[38;2;252;238;238miZgqqqqqqEB \033[38;2;252;172;172m.vrrrrrrrrrrrrrrrrrrrrrrrrrrr777vv7i.  \033[38;2;252;238;238m :PBBBBPqqqEQ\033[38;2;252;172;172miir77:  \033[38;2;252;238;238m:BB:  .rBPqqEBB. iBZB. Rr        ");
$display("\033[38;2;252;238;238m                    iM.:\033[38;2;252;172;172mv7rrrrrrrri\033[38;2;252;238;238mUQPqqqqqPBi\033[38;2;252;172;172m i7rrrrrrrrrrrrrrrrrrrrrrrrr77777i.   \033[38;2;252;238;238m.  :BddPqqqqEg\033[38;2;252;172;172miir7. \033[38;2;252;238;238mrBBPqBBP. :BXKqgB  BBB. 2r         ");
$display("\033[38;2;252;238;238m                     :U:.\033[38;2;252;172;172miv77rrrrri\033[38;2;252;238;238mrBPqqqqqqPB: \033[38;2;252;172;172m:7777rrrrrrrrrrrrrrr777777ri.   \033[38;2;252;238;238m.:uBBBBZPqqqqqqPQL\033[38;2;252;172;172mirr77 \033[38;2;252;238;238m.BZqqPB:  qMqqPB. Yv:  Ur          ");
$display("\033[38;2;252;238;238m                       1L:.\033[38;2;252;172;172m:77v77rii\033[38;2;252;238;238mqQPqqqqqPbBi \033[38;2;252;172;172m .ir777777777777777ri:..   \033[38;2;252;238;238m.:rBBBRPPPPPqqqqqqqgQ\033[38;2;252;172;172miirr7vr \033[38;2;252;238;238m:BqXQ: .BQPZBBq ...:vv.           ");
$display("\033[38;2;252;238;238m                         LJi..\033[38;2;252;172;172m::r7rii\033[38;2;252;238;238mRgKPPPPqPqBB:.  \033[38;2;252;172;172m ............     \033[38;2;252;238;238m..:rBBBBPPqqKKKKqqqPPqPbB1\033[38;2;252;172;172mrvvvvvr  \033[38;2;252;238;238mBEEDQBBBBBRri. 7JLi              ");
$display("\033[38;2;252;238;238m                           .jL\033[38;2;252;172;172m  777rrr\033[38;2;252;238;238mBBBBBBgEPPEBBBvri:::::::::irrrbBBBBBBDPPPPqqqqqqXPPZQBBBBr\033[38;2;252;172;172m.......\033[38;2;252;238;238m.:BBBBg1ri:....:rIr                 ");
$display("\033[38;2;252;238;238m                            vI \033[38;2;252;172;172m:irrr:....\033[38;2;252;238;238m:rrEBBBBBBBBBBBBBBBBBBBBBBBBBBBBBQQBBBBBBBBBBBBBQr\033[38;2;252;172;172mi:...:.   \033[38;2;252;238;238m.:ii:.. .:.:irri::                    ");
$display("\033[38;2;252;238;238m                             71vi\033[38;2;252;172;172m:::irrr::....\033[38;2;252;238;238m    ...:..::::irrr7777777777777rrii::....  ..::irvrr7sUJYv7777v7ii..                         ");
$display("\033[38;2;252;238;238m                               .i777i. ..:rrri77rriiiiiii:::::::...............:::iiirr7vrrr:.                                             ");
$display("\033[38;2;252;238;238m                                                      .::::::::::::::::::::::::::::::                                                      \033[m");
end endtask

endmodule
