//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
grkA0BvEUO/TYN+idVNmaoNxCgrdqsM4cYVC5fg07S9mwx/rm/n7Rd5e3enZXE2Z
AHh7LrtwxPMXtJebaxU76HbG5j6COBvDRmCCnen2lzzylu77NCeiEOSBRVCssOpx
et2usAGJnwmbcTtQBjR93lolfoKiFGMUdRCj5alx4g8k+PEM+uLii+vPlivNgays
WNMUQ/8S/Z4M1TmdT89wB7BOXXL2A7kQYljmNPy8Xjp6E0MKqv+tDx/ROBuTfxgV
U4TG2HLeyXkqYzaR4z4HawSgC1IUvMWj/kyyi5B8iLp4AvP/sEKKdu1aK1Ii9cEZ
82zWN499LoI0ZJVJh4Yp/w==
//pragma protect end_key_block
//pragma protect digest_block
PHOwabowR1VADy1BltHB3Dbl6WM=
//pragma protect end_digest_block
//pragma protect data_block
NfiOASyl+X99QbALW9Vq41oQ/0HD9oA+wFgtdf2KH7U0TXNLTVgt0jvfMZkj+T11
vUo/9VKo6GXl7ravt2dByBiaJf4KQDAxnCD7Rdk7T4y6Meji7DrEsjybt4QxuQU7
mOQI3TIe6xrR1PScD3zPgbBqU/+kPr4ysE2NMj9h8WvWP1xIjL93hxrHLEC4nuN8
QxjwFsHYmK8pwVCZx+By82q+UNZ2pehK29SMRMERMh9c/D0Ifxb5dKBSdiW7fi/c
dhkzn2B2xioiFTksYoUSZIFWNEP7b4YmoIf4w3smgbTRtsNHoRuGOgP2E9b2QpeO
Jkk9IzEJByQokx7i2LZuovWcUUBH5pYd+mSgbRvUIN2jOjqf2sZzl+hFzS+h74pY
66VeImPZZrjGfVpCh4CP80IvZfVq8sHQ4CqnCkf5KBTorjZAY1uTcLLeb0lYuuDK
71uAhMJBaXAckrQhydgxxTn7sYvkK/nCkJyqLhnU+jcvzozft3L+zKhhQm2ts5NK
l/+EOuRnvQAPVdkW5EhWulYIHFSctmmKq7sku4oE5HJd/K1OL9ITWeCYbD3IeHwA
tucIPHIsM8PbeXKyTCTh5OUJWttcA4PbK0JCDu2enqvd2MqEpdx6duDOZCAnZMyC
P5eCY5qTvdAVZCNRMOZHM0dw9h/CetvvEEL3L4BDCG4C8zM1mtbodM/OvixsIPvx
ZZlH8L1dWJn5xlsuq04wbsnsnySWPGpwi3sleAYlyqRsoMk3dFVqnOVaLtIVTB5L
8D+gZA5jtW9DQPd8C4MPu7L5zfzroqp1WpZ3Pjn9D3stmuyPUJPAL5BAn9TEeIFk
pK61rLGIrcWJPQuT7YuYu4bZ6iTL3hJ/7nlPPkkhbC8c4pqOVtXVRh9AKG8W3Y+1
nNiZ8VFX15EoR8kIvB2Nr1A6HFR1sBiQkVZ51cxTWd2/2vOxbB6P9VZCcNwVWX1+
fe9R8LGTWV1YXjIL3lX7OnK5jApA8wtWmgJ473IEpk1DLefvC6+jkefTm6vfJMpf
fXfBbIafqDbOBf0EKjmobXizQEDejmIF16UTSECndOq9FBskmAk5RE5mYWDgzdQ7
668AsrRKllX4kNKCh/9cRZokeBrdpps/sBYUIsa9FlKA4D8KLIyTMGS8f/cqWjsV
XtIB2DDizvXlXuLOqXPCnU4QbiwalxZmSPgQT0toDl9HpTtqsd0bbtuLpCRJELyk
qd9Me0qDl0pA68lhB+XOLoj/4/DiC1la7uzlsFoB3jq7Hs4QM/MYEXygQD4LARde
Qw9uZTUfMy4gC0DjEIGlFhHO3KKPkOoH1PfAGeaL7lK2FjHKak+RNy7SdUGMXh9Z
X/cQ11kQozdT48wleXFvI+e8Iei6GBLvwaV4lOdGBMQGLEAtks3NBnh8i2MyCxF/
4BIlI+LgFI+Uu+CZ4V5sBUR00YcVBygY7XFbvlpjJeQ4GNK5rOxosCZtXAhbWGzp
0dtX7euVCjYjJkDLLRJ3gIVRibvpgiwc4gElNr6+GxOsMWVpQRarjQlz5Lz6u1JL
huoU5Eqv68cWvn/b2K6f4D0FS0onuPfoacpFaPl8h0A4YpFv7aLSZuqTK8Jh9LHB
Xzw1KlvICBDipD5LZpM2ocC6MvfV7dwNwccW2oVK5k2Mr78oWsqEPS2cKhlE7Mfa
IQKNe7POFjxPszkoyklmJnAkxfzUZcWp4UloCb0IrEfNUAoAmOkHDEjVZbmbWlDV
qojrK4nVhhsdCiVUvBzQIsBl/hvvTN5vnKOWxgn6eCd9TEGymsnD728oUxTzpIZU
WKkQP0Zp1LoYG944qFzajF/Tti1zqiKtgR5EFh6Y5V/kqzm6xfmm69ZpyoyuatOX
0DDqUJ3kaI9RBmdXOCcNWWee+4N5ttF1lBW6M58NGc5k1o3jzqiBbVouu4Qo3/Ce
UneJtiNsfJ6TCilwXbuvvJDaI/2USoS1gHQgab5ZncJSC4y281gF3eQYOGxjqFUc
1fIPMQp/3Ck52A7hWzZ12uhn465jyeWM9Qp06LBHdPPvp1DrVs3lU2YWKJnaCliI
NFUUdQjFcKO0SnKZISZA9wF9R9g/B3bJ/fM109XrBcFFJRYuPt+pYoTiiE0l0SoD
dT97alvVzs9gH4fQp1JX4TCKhA0dhMMYfaTOpv49oY9H+Czo1tc0yE4G793LnzHK
b9OHCvpVnO20Pw+yyfeJbBGxo16f7XLb0VvU/LWI2cPKryDIlQEiHrpYGS/JuXiG
+1V08M4VKEQfuNXYERz5BsToe0Ej7ZQjOyOCD/P8LxWLi/TKI0fVcBzdFACO76zm
UuezQ7hzMVP78DC6siRB66jg+TtU3JJt8PdOfbk69VyVRdMiV1V/ts/Vq8olXbxN
3Rp48sERD8jUWbN5qVK5+XaoSFIQGGSSdIix7xPjKH7VUI8WojiydRCjeGYPffBw
DkWIaCbulYUfQoVD/31Uf9D08HpBxJYxRjUWo7WUf1Mhlu7Ml34tmjIlfgJ2LPsn
ZrpbFRLGHBeCuZzYmsjtWKi0XW6qjcvIETG/qh7w3QmXjo56hzvkE4Yj7Ax6Qtkh
Z+iyvpa+9zGspuPF3uQ4IKcw57LyZjUkxLENv/izNV5ZFsEDCkP0eq9I5pEzzt0i
EYrei96KdZWrgmPK+R77+V4+Ya5FHwoPtfVZG2DQcFOQsfpR2Qtgw+9HUCdhXogn
mhy/uQV//HLsQk/Ett3z3QbmYGYcrsQ8VE6d70nuXaoJf5AsT958BkIuCEuGzo1g
L2e9IhslagelxdLYz+J+fjIuSxuHAH0v6X9OnBFabcfwpk7qBMKHtOYryM5z5Gdh
/Q60ixdY82t4hIXw1e6UEQ794k06jbEVsj4HuosKhUIaw/Q62iBmUrUg0JeL9lCC
0wobC+S85DoUrqSxRBNtsnnqnTyFMwnll54xHvmq2+O2THRoUMXWnyJu7r3hgsxP
uI7ctGdARr6aY99jd4RVvcgr3IUAlIZTtmYgyMAU2h6+TtxouZCVSQIWhyPQ+zZ/
8MnQfu/J4DtBTiXmWMo/ZLQNXhFKykhKZVPuY9loZnuXmBBmCIkyh/JzG8p3g1F+
+q5TyOXOhJffq68BBsGOQasWprTlDE0B8qsFmVS+cbALmzDuau+apojFg8ZRgLYP
6zOMMjRKc2TkQQndSGfk1UDz414MnRHfxjONfg2fMz+rRDhRsDkhT7+MtXhVdy11
15s3vHfkMPDObJM21iq7PbPuoR3c2DK2hfpLJ2kb6lWRbFR98tJuLv8bA5cyTfLm
CBtsfX9AG/RXnECHjXtOhTDgiJzUzMmk6A44zaSng5XREwy0Uc+NXlwobO/vZaRv
5CIqspnDcsCzcsd3+CLLkkBKNLANJXAa2XaGlvBLl+uEVOgUbcyM8nUvb+Vvrot2
gZ8fhtL4Ym1wE44nveC974iQN6z51zURHpCv7VJuAJlI6o3EMCXgcmoJVzmg7fpW
bfo3RQU1CaXEk5BmkG2WqOhQoZ2A0brurKQegp96PcoFXDMgqtuBOhnxgafS+XNM
SlJu2NMSYAYlCHq4CR3UVc+6LR3GLrq2kG1yAuBmuG7g3gTOegTgcjoDNj0spYi/
ChJx253MqiB8uDWW6z9+p3skfGxke9Vya2veyx8qmfJJjWyKF6Cs/YtwoHyjiYp8
YzHg669g61dOFxZ0reu7EjCec2OUiM/C+rf9CKGBLQ2Mwqzk9IBALm3XKWN5jFBz
wwBE6vtDSI37P+MYoGHwLskbTGkh0KNxnt/MIZNvEjj6bgIzhGFTwlr4r4p1OVSF
Sv6CQMbpgl94/nroGIEGfyjejHRu+i8N2gmZG360VBe10zmdX3aqyUZHbimMMOqg
uCdLw5UY4pK1addAtT8YdjzDqHKGAtbVKjjE4dg8dULvQ0xHcGgBS5s4Q68JHk1W
1cwjX6PlTPzVLHEr11ikV3hao1FLbduR5uXyVYaRTnXR32KGW3OdYJ0EkBLRHfWJ
O3+r7jGgz15hUi3UAjZb2hWdBb/bBjXa7dVhPBlDzSQnCtUnthtB7bIKXdAXHc16
leRvqT+4QXJIoo96TZA5KZYKwBwQp9yyxdK/SEZlHUXM/Bt7pcuc7a9eS6AgeH/6
XSfzHnWaZJTjr5nDDlWJ4WoI1tSMfIHGDMDc+k6F/TbSOqe6aUVabAcBURvX7Mm/
ArJh1CLMbhrzzN/ruF7NEhUmnhGYu31j22I9PN1yotifjtNbN+utEPvWvqXS0rNZ
+bn84NbNjrdx2x3yFbxr8nh2cE1mvDGkGgsNUg0Jwh/L8wMnPniMi0HEAV1Uu4Xy
+lYnGm3LTJ1b6y3zP50846xsWK5l/+votVx5DLcpJq/ADBj0IQdcdEy8uY4SvwtP
uPMKi71ZAzga9gm0eTJxj87mubOGEQAj8xVRH5efFa9SPkaw3OmqdCrUldE5v+Gt
xlg77k27itB34N3SW76nK12DqXW+b2CbF77Qka2qO6f/mGlalA/HEJh1E723zsJs
pjYLgZWuRDzYJcGK3p6pNtbwayN8zIYH8QuUgAjg7YFvNYe9l6NXBuQ/bK1u6a3Q
Q5BhegVdPG7DuaqyAx+pneJs2LkpQHJnhQ57l3Gb7FF5XgKM3fa3Qiz1oh4zN23R
DEfy6JUZ5IUKs3pplxhJuFi3qxpD4dk7eBfnrN+hwkfDDn5VOJJqd4jsjHxTUAyI
c9EBa+8FN1SM4anDagL8YcJdTailStcxGVD0+LBRmbf0zntdMKaZ+eQynWByQqZw
Ja3sPy2qTAhv2WkEcltgbXAIUxzVV+CyUxHUVTcXLqau2Sj34A0xMPR6OFf/kZw4
FgBVoV4vufAPqWulp62O8pJDiJGY0cCVGO5sQS9i0+LBSuCXUWN22AUgoFYH8cWr
pXsG11CSzMf1WYv0n4ZnCn6KFa6I+jEnRxeQZdF/xr76N6Cm5Eya34kEMwtXk/l0
BRdEHArYqeOr3Y/Kgx4YI6uYokozszHUaRG08KC05wv0gzAYv174xZ54NbOGGag/
k4kPAjC4xda7U6AW+VW+lGVbrc1uFWKAo1CeIYFciZ7/O6Lqg2CCtHEoZwhSndIs
n4lgdeOOYZtbs9DDVI2Lh1k778AjCWyJsT9SRTrV/M+9VQZHW44rjQqX6ywySVzQ
XKEHnCTEQbELW4dOAqSkzTnoKRlXVsmUlPXLQmBIye0CJcdNxUr/5BjpzrO9LGeh
GeODmMlhdacne4B4KJL+NQYrEU1cmWq3CoT0lzS84uzoYRA+qR+t6e2p/QKfHp5S
b+Yklp92x/g7FzDXnu0iDJt8pBCTYrBzrDoC4Ve83ClyTkGuuUd/H7dYd1WH5QGW
us16O2rnfQLB7S9tTgMdfNcHq0cbRZfpTCPXYp/TamCqghx1eOSgWEIrQzaKwfoq
Tehze+NNgmrpcH3JVCY9QwqlW8b/uJGe/4WSTPcJXpgfSNmdMl8ty14nEjAj6PR6
HIcxqbMXtoIE0bX8jLwa/0auJhwFN6Bw/X7XCzAKxESa0lbZY0ghwRWNxcp9kKTV
LlvNqt0K8Uyvs+4ZU8etXzbwa1wmLN9TIC5UTAx1+9/xMe5sLrI5ZCT9V1xl42VL
mTyGGTu2z2ooefE2T/Ouojyukc37Zivm3puC+B+FBtFRbWV45hiRKrSXYBx556gS
1hpCYSp/VGBW2Ga66qXFh3b//MIRFzbl+Zb4LJg3qdFT+AdSMRGBM2mf6s1r7n3j
mecfHDqh3YsjH6WX1BumgkjY6/fCmAf8CBNWx+hIC1j98HmoL/u16vEVvT6G2J7T
dkcqAgMG3/dwWwE2IEh2TxRqCSzmwVQhKjLFcJJ53f6GeiP7Egr5H44xczg7vDtD
sr5cq81C58sCuy8pQA8RViMhYgYpXma8hgMA/BuNdpmypoD1RYxaN2eELkL6zlj7
0Tps39XeuUJ7COBethDsNFRU2e2t/AoCMZ24mknKGWsfWZd8o/3Dk+9t893EP0eS
xEivcNEWdYtsxes2YLqPl0MwVrAaLAaq9O7ehjYA2nWG78Nx3X6cqYCIBBQTFPZa
yxktqe1ZzezamcArOGyj1CpxncdkrogCjJ5gM4SzjB0vC8LanizbaW5cMbWGDWBk
8jO10BQdUbB7VwKrb3MddafGaFCR8d4STrh/D7dBYVazU8VwqBAKf9WPF1jzzUko
K03zeuM8tfss4WJdadQ8E32yNGwIwBXVc8O10i7RQ3FjqFF6mfMQQ3ejV+Tn8HJa
moGS0d/U93gHSeUmSP1/PxVhtyoyEomSHN/DB3bOoygVmWoTFyF0K3+ekNOXdXph
uIUzwfrkMhVQb1VCAOU7dHInwl2R9m+/fPLE9muwI6kFgr94uQYtfl+RnEri28WQ
6drivWEVDMDzy2dTW+hLVZ143X709rGYEm+qlJzdOF8eHQudlHQovXfheIX0Y7Gx
VQnYDvZLva4T7B3BruznmDUTwCa2/NZbE0CT2wyzADRGIyOfoTlCWsnsRhWq85+9
NttI6wNln3p92WPjHhexvZ05oGeg1MuB7b7zg2rEI5FNfoS0J6jiPfp7/b7ch9Lt
YaE3oMmIhgfhtIZoM9QFZBjp+k7sGsLfAEBYjbaMYwPDFTmxLU93u0ty351/KaXY
DbPnupCOR6ELMz/Je7tJk1m7qLg7nnBwM0quANzWLdzrv4Mdfk7B9fLz1BIkEsYx
Q4wdg/JSf7fF1Wi4CHUa3SIPw50V1vK5CDKhfIkl3EkFi9ebD8lhI5Cxz6XU7NDH
/N3tKP6BJ+lBrBerPrtVISr5+p2Kc4fWwRfKG9GgVsFfJ6Cpw/5mHTrcdrftrMyL
9YvosrOGurGu5liUd2QAQvsI+MlpKKwJIVqATM2AMf91/L5Xi9RFmWD4vH4FsOXL
07J4RT5okFVy7HkQAMfW4y2DIuM/5hNWKFUy9dY7WkIqdcEWBjAsLlWLv7S/+czv
nc9+tVKaVOaw0ISqAPY+GgQEEMBH1wDvAdeG42I7gRvQ+2++lomJDJbLqM4TTAuh
7pCB4KkAHfVlhs/HjQe5Sd/q8zDkVjKwbVCVm+CN/3UIDCr9+NXvlRD4k5I7STZE
lTNSPMtTm8zjfypYS0XxQEODDkHfHx5QPAjezmlZHRNteb06PMDzsA0KdguQA7o6
RrZiF2vxkeTKvJq+OAwRKXNfUdvvhJ59tilQu23BKVvGFi/1FoArtmIjLR2fDl5k
IRym7qt+0M6e1SzqPqsQXOOGb0q2j7g2htHUDPMT7bQjloJj0R9jBYz8pXFAaFXk
O8fEs/5P6pFVgY/8aLq3U1HJq0Xof8tJbTIXAPqLO4fwfwiT8jfHsTE7B44XwWs8
2n8qqz8+jei9L/7U9a99MHXHvrVrw8w6HEKu1nXFDhN12bHaNGcm/feeZ5o5Ermq
Mtcu4HxBBceMDDbaF3375X5DAmTVU4hONt5H2oAb0Sfa554QGi+fMgYGD9VMgm9/
NzIRBDK2fIlCwdVylK690O5JT60SZAkJAVi4bWG93KN/RSa590xE27SaDxs48B1f
gjHrlZXEQ4fC+MrD59tsAFOYRdSQEBdH8isOVSD1c8p9FeOx65Cfg+XDvcYrN4Y6
8GDbbk8HJ7RB6cMwCmrQSCD8QNfDaryu7sBr6Kmm9gCXDMbVWW8edzXYK0sT2Ndg
LMXoWAcxL4Noo0ni82mQsQzn6hB4no6p+I41Yog3SEMrWB9tKLk+sz1tQJvK7OxD
79smH/ptQHeCq2zNuVt6GV2rCS6ZpshjdE/4X9geWjkOCl3mPSSHwPo/c5xGfWjH
GnndSGQQbhkf2+1ga6ei+hMOc6VKr98VfBrqGnZ7tAlLslyr7zMY4TdMfjmFSxzA
X8Lxb2HjJf5P9mpETCUU7zDgQmrgePtPb8jmiq/4/Fe4jOyi34Q4NQZGW8ZU3k53
cbGIyCWkINr1qSEaRirGubgL9Nbq8aDkHCIxurjhvtJzn782V+pEhXLkEUJ73HJv
fs9AnaJZY5m7MmdQHC0oaxDXrV03OehdtlAfQ14iwikKqchoH873LAZy2gw+eSyA
MjXmwL3Mpil1Fctb6GMEwrj6wirx0dWoE+UZwR1kF1KYr5ouNnVlGdCeqtn/WOvg
OT2qA++NjIACxy5V179o0xaVH2fGNaUs4d2cFC/KPzTXOh9Hx5wvR4zvtK/2L15s
VXMrY7H/2qpXqd/i2PNmqZkQxjRoA8BMvmkS/dGTC1s9GHH9r19oXindA+vjjBcP
oWkTNLSU/1u2uxR0zB3eosANq7wcvlhI4BqglHTMz6p1gHftJzQq6nuand5OW+np
zmnskw5r8yFxMuy6Ug4WAJCN5mlu+dD8NWD3jX3B9CIyAVntE6wYv8Vcoou4lxix
67oJA4hqskqoLQNMSru0OYUD0iOMjcdqv2QSVa2iwxvYLuXH8CRni2eKjET1uqIW
qcme7T+AnJHnTYO7W5XJ0RVCojoQiUtxYGaIWlj/B4wLNHagyFk9k9sTtPeygQ8S
ua5cxr6Z5wAzWD8VZmXDm/pWm8vPfyMRVq6pglA5YM7T4m/nfhS1LQNedTds10Uk
+Nt3o7QmifDAiJLOr0YXkB60Q1w6EbNZkwl2lp1Dsg57iVbj22Hdr+SegkU+QaC7
tY83eHoOwhSzraCQGAImAUwG1JdraY5iZtxXhq9mYChe/3i/MWW1CswZOy9ZrRCL
+SASZKvBP8zHfhCWWqzoVzTStFPwTSuHUzwEtRSqk89g8IhqEYmG4aIqWkjehryf
KnMVUMtRxVFsjt7NnrP+uc1/lIjGThS9HGuKOcjAX7H0st/oehaP4F2Og5Is3Do4
hDsQU/9TrVE5m6hn2zo5aGCfXYxLCmk81pzzzfyqPnqSaeyhiS4428XciTDw1E0c
lbr47tO+0gCpxs1w4ccWu8A5bq2lIOsoxrH7vAMXnheogvePQ+GWgVpjKwKEKyr5
/Kx+KECoDM9A2daOjM+HgGMudzdS+IaH3xnXx6EaGMx0ePM+kXOIWnPVbiIh/xgT
/c6IzzofRob6SRpo/QXysDusEzoz8npbpKTzjIxxLPKYdpTQ4rNGPOyWwtGTEYRS
l8lI4O95fX4+RMoNt6WT+03ne44egXDZigABajjCVkhY62CCdJQwwVOpYVz4zoiJ
vV1N4Z4lFrRw2YymXKfmj3d/AB1vD8I2YUrBMh19GlN6JNDxSEzBUs/lbhG5HKVD
aCypuXf7VLWJu25lWp3fc8Ha9kpVGTRIqiFSlIVP64rRuRzNz4sHkB/jTIzIt2t4
wBkqAxzAcfkkXbnu3mNotHJqxBYa1z7iOjn6NJ0nzb+0gc5NtCosm2MAsTjzwT5T
uid5Q2Jj+nvKxyXIzxGth2uqIbi9giEfJ+t12FGeT63dkNa1TEAcdBNN2GWC+BBK
1kr+iXse+Nt4SzVJPtnQaQ9XwJ6A3gY0gtkpehY2iSa9bW/KMHp1GylQ9E8tILw8
xku0Ruesn1XtTyyqvdc9r04c0Uxr3mffq0sUaYkKhA+1JtmLO2BdZ+I7eoJ1v5SF
cNL0CbSbGxwAJDXaVfvnVDWrauQ1JVW6BTd2tha7LeW+cb/doP2TJ7eKF4MnHove
O48g+FkUeZCnvUMcdsOPmah4pWDEFErt24rr7kGXX2FA9b5bsWl6Xvgjx5ZRNumh
HsbeKym1g+dM8pv97wzx1jWqH2IgcvUJF62hQ7I02aTLPXMi2Cz4dyAjMRES3y1p
3hxDp8jkYI5kkKzUchKb2wIiienNfWFqThgIIU62W/tHtkPoLlPAK4IyyE/5iM3k
TKpKQ0qv80IIcwsgxP7VUqKKIAhExEs0maktkyCZasljJZYd01fZLf7Vip1YGMJ7
WmHxoSUXJ6qMObLQGf0VKQmHN42P5pbonuNTZQ3jHKdssgZhl4YGrM2UIh9UO40a
msrsQJe5RLFIzWiWrz3FI70/ZnrB/jj5rEGXo7LSdAJf7cuj6T4WYJD/+Umk6Abv
cjjYb30sLRdKwZnpq5QpJaT0XZqv1TJpdDVEqqwPR1qkxONFv/rzBNi/Q4LY86xV
kyp36+Xpi4ibt2F3mpl0qKh0XB730aNP01ojWDS2jpcUieEYLPM2Xa0UoV05gS/6
s2Zub6qX4wemSYAERiMGhZmbgN5FTYk3A/HjzQG6/WdcNTQ9cRCGvd4uoEO6kklz
noTtXXKDetS6rYqy0LSYn+kfXWpjGv8GJomL1U/USxsbm1LdqYBNFEIqdKic/pZx
MWwG2ESukxV3778scBVWI8KVUI3GIg1gcoGD32xvS4D/VkvVhThMnowQ0TuCiQt4
EG6IA2nAj1jbjBbUNEVkPubzfqc0cQ3Ql7w4rkvWa++P6DWMWHndPQNyKAArmubx
+tSAXUHLEMEVJFHnXShYky7FOfqvcfK0YvC9OwkwWWcXwrEGgV8KxnVvR4sMZ07m
Fm/CA0Yh3rsxLTF6YqGAQlxc2ZLYNNOd2dJqcBgNQdDsxd3Wz+yHiWER7dqYVDSm
f6bjp6JPw4BDmP2YvWPBHrj/AWqir2jcHEJN1VSukB5U8C9ZXS+K+4xpUG98xk3D
E7G3OjsDO8f6L6kdAUfweKZb4qGoJhek5SQOhSC4AQzpiBmne0Bk9pDQ+Wg6Ob/X
AePUl+oTS3LJyrVSkrloYnSy+fx8geYhpdQr+CU6IfNEZ0MBKLvbjhCdGwHJOS5+
2YgvFdvvuAMTfXHuzWfoAViFWRFeIw9Y4he2EOUz43+X46fGNgefchQu5gR+3D+/
fN+Tvm/Y06QrlbB1liEgYE2BmB3TLSOZ/axTqrZvSEl3yDbu2FmX3+j99j9aK3Lc
Ib/fpxXn7J1lN2SoamArSaRYEgvH/QQlOZOJugBIxBLwFoZS5sliGLPapjTIiiv8
AA60dip1X6yyHotBEvZ7RxLTk2gir9ZabmKfcdTopr27gxGTmNB/LFiglhsHhH1x
sDKhd5YQjoFW0jqIp1jVgNYrB1LKSyrhqb9YG+3zinXBZyOb81v+f8u0/eUe0WW5
EcXFz9Vxpamq59A8vJA64qWnaEzTDkA/9Qup5xtQmry9wbAilx6gjhRQUPCJ+Qeu
SBzflTEbxuiuCjndxrp/YPMJhhGrLEL5GvYEFfWHmYCfyDjyGaHAuO0xm6umahah
HN5w91wggUTFE3UGetfFrRZ7qSwW86ScTZBXUR5E+rrpXdhjwFBc+kTauvT4AjKW
PQDBFPdt21LphVHmRQsir9NTx0ORRwgWsaq1IovHL9ZMqgA3COvqUcKjH7BrmnYh
ZjTkYO4TiYgUPJQ0DN9dc2bLAAkxStHajI75tQgwZmCRCUANw5sd6+EP8nMlyAQv
dYFhKZ+HUxyzq4awdB7/D4uA3+y8Fj60KFrLARuZdO4wNarTt7gvzz+7ybdUUYll
KtHycpCmEOUbmejak/tQj6Hp+Pf4rJ2mKpBxPR9j06sxp1j3GoKyTnyujli7Pn2O
oE75wBoSdWk3cFYJggpY/JoBOEjGWhucIh7kL+DezoxqGUxmhqI+yceHhZENeCis
+MAxuxiTisMGLOmi+tpPbymlmV4RbtXg0JMQPfTwjz8X89dOLJ8KFqraX/lIDnV6
4sAib1QiN9s6CmPdGd6Gq/XHE/tuNXwn88io/NXQ9HdX1ZM6RVTbSgvsCRm6vW48
zE8krJehKHmaASju7vZpxqvZakKg5ihI8MriAh3m3cBbLubWkeafZY15hsC96Nra
WsEmdTaEll0sgV65js0XqhFY/zntWiyjIIldaZXhYTCyFfdvZIS3ulB1ySRWh0H2
PE6fPxQunXXEU68aRfd03Ytx+eRHT7Xx8Xl9W2Q8CrS64rIWM1q27DgD4pZMhyMN
2nyN0Wo7PlqD9p4kegJUUmA6V30oJBJd5a/+jRCTTrBu0XDAAUie97E1A+zkb3ui
zobuVPwUVHOToN+DbjMz31Hg0v86AbfFcyC8swj5auC2rhUqRIpQqoLU3ODKQbAn
/zfpSbOTyD4PB4xyCPrP8S8Oovb8URYcJD/ccjT0VxmoQ+pmBDMYGiyvsE25opz2
NmYIhHZaBHHjRzLz7HzLCfTopv5zzoNtFzv2mFpaULbZoWvkukjQjRZS42Sreo94
Rmo0aQ6F6vL3I+/SGA/2rJVdsY7zNRgjUgg4fGPNNHDFkFDMdhz71/RlVEuczKCg
iokYpVpqpINq+mCF26pEfs//4mjBsaZ6scLajEfzY7hcLZWdtI1pEuA27tFqcDOT
T+CX//EWKHF/lEqbeHfLgNRcdlmQ2sHv7lQfn4PP5yjf7t4O4VGo+EcmDScmXhnG
htwZHun5nYC4Y2b3qzpp4qHOk0eIysHcfhSCxjovS080Bd/rDRtXTFJZP+0H/MRo
EzYCnQUuyMpOa3tcVMdC80PIDiTrigIUcblPTRQ7GFn6MDFzGdW0eMX7pEnwc502
TTtH9I/8eHyeCv9CrId/CdfstgfEl0oYk4kD02XPcqO68KV59DVQ54lOn9BKiiHK
yfo4jnTtcgr1qYD22eRvoU+pSAWLN8fioiRKl7o6A8WAzciId9ESBMOcfDDmZdOW
C5rmR0bg5C0eHaF5svRudYpGvZYEcf47zadqmdmA3zH32xb1I13BnGOuZL6ZTIiX
MrClSSCPMLcWXxHXczYekBDrl1aBd21spNWou5vKYIUnTS0CuvytJsUWt5cIgEjc
wYo6qodlNtekRRGGpm5oiMEaJc7E/mpIZ0cYUp8e3qP5qpDRZsMZqhLlUn9necbR
058tGK8H9m7Ap4xh2kbE1+zKxyCvt8w65Chi/Otr7x0QBCciYiozGja8r9SILWsG
RbAcLSzCLOOfk9ye8UATtXxdyAFfYbI5lRrXZn8h0oh5Qx4jYV24DZ0fDrEDDJye
JIr9NYVzsRh4pms2+kAowjiswHXAX0dRRmO5fFsQVO9B9v9LKKsTAHjhE0ATHen9
rp5eCbw5IiLQSE3PqHJPleH5GUS9ajsAIRasKnmmVM3QpMe0EYn0uXDlLP6bPHXl
ix0yDUjYGH2xwV/YHqYPqSLJAWCtlCi5PERY67oaxuhXrIQk4oHX9MKDQO0RntSJ
vp3hpj6tQkF6BThSbp4MWhwPI0d3E4bFavRAkITs81Pbo/ZF+BPjDw2B5UYxzaXF
c/M3XQ5CoecWUEzlh8f1HZpl6ec/xLLYlqDMiCqkFbAoKWkYMUgBzwPhAZk8ynMi
6NudkovKxx/JCPjrQoKnK4Elcp6ldHJZ48ew5DwCKkONuOIF4o7wKdWnTH8qexbO
dBmgfiMvaUUDMspGvEgEa/j2Rlxw1CrsKu+JZgHDKIf4bKQnixO61lZPe6A3zhvt
WlOfv5VxRzq2Npr+Tbv5Knp/fPnx28c3W+uPKY83rqwRDCmkjwMrQq8UDl6SASI2
RsknSaodGbSqVE3j0tkP2YijcDQ6j6j8VyPZPCssqk3NI2X25Q/bNz+LDKdRDa7/
etIYfrmyLFYh8UTwmyfBPifS4n/Rs7d4tGCNKLJsVmRpHFUa96vsfOTmdf/QIdQq
Ys0Zg/FXffIjc5VMQKkKQuVuVJrzUWbOnV2nMSJT1z7wtOsGIuLUTuX5WFFZuqAp
VlZsxJVCSpw80OOsp4iT/1qZIeelp81tKiO/vg+2KFo8MrgdJCMteEeyfxsFSCgz
/4q24e9hrDms0ksbYBq+KTPNV+FWaMLVdTftDGsg30demLlfx42Kqg6j8dBW8sbC
vqgeGTQVf/hpTEC36DAELzHG8j277gik+Tua0NnBpXB6zTsEK5xX//a6knGo9quD
4RFy9b+b9ln/ptdRqOd2aLtcZ+CJNwLEpIL7IeZ1JAV+7Iuk0JcmDU9xDx2JEWDQ
a6j0uR27CRz3n1z3dlxUP5lV5lbtXFMoMS2KaZZHr+6T29rYjqm7pqs2YYTivgNd
DClzXCslc5+UosJkMEd6NpJMZYFrV/IAfFg1THTiABCz6Fko1KhusMxdelpg+Lt1
TnTQZlUSxk04E5dDONlzOwb/cQgyUR4uTNqsdYR1eFG/nWoq5DJtzIfHzxT49mcS
URXgZUbL2DFV2SviQ+OEuXYB0Iud6tT/0PNVEpVHniIZeL02qBvXUfNkuwODZ9SH
zfy6nHfbnuKq0xPxGoqXR+1qJWKOxSzG5nrMJ8ArTS3RrJSihjqq5m+JdRCACYIV
nuoHlSN5A/GFw6uDtTD6wMQC/WRFT4EwbfcfBVhtJ2CvstnCaSnjWpD93UOecutA
ot5OCsQjCvEbImgPowWKR94J9wmQpV9GqId554PHreKni5VpBYMENK3GE6TUbTp4
jtZfUVNSgt7ME2c/8UR0ESrpDFqGoKPsotSbR0ix7VynGYGuJ055kgI3D5m02qoJ
TGa/kPJdhMR39YVl3hAouZKnXWXpjVOsqC6Pv7QqJzpD3hwXvCJFPDeemLuHuq2J
LylKGIyTfKfAJQ6NKibE3FV3KrqmgRFAUXQoeFpFdyJcW0biQ+F6q/GfJL+MxfX0
ed598qCQqrpGADAiyfFsunIuIlLNlVMf00Y/r/wYCx+3f6MEK54oz8+dj5PN/EU7
Q0vv7oWZ6/zh2kS8bNqmlWMAox0Uta/RwU1Tv8gyYia9Mhjr6+7exOcE3t9MGzVZ
ZeGUhutSOvtAWDsdURL1QqC0LSgwODbg7oCDzwUkDY3/SgcPW6+UPGltuRpasvYK
uWIcDkoeJBcnXwd4t8wFmPj93pBx62dGlLrVBMT7MP294Cu0Fnfhv9SVHE9ZDlwz
+AENsKuL/wSVLnRgHPxCKBjv1prqGcJchs84fdGmUwKkWupAc/52oezFZJf8bTfO
R5ocU8AAaW0ObOnp+QxDR0qdbGTTKXghnSW0jy/o4VjHXtnVuwQ0h/vIuJBHamGT
QonYJIfk7rP5pfOceY2RpS+MIMhEWPbvDk7ITXRK8h1/HH5z0W9dT5+Z0Eg+Bfm3
5G4PmTJnwUwkyNCc7BbGr79t/X5BEaX3TWAQCIUcYRiKAPP22LuONXimG5IvtuzF
Gay+ThI+a7jFOjDHU33aLEi0cyFKPPSE24iRcRUNmjAOTGG4Wj4soE48ZVdTzGxe
mD95m37TC9R7Sds0NwjNEAKJXtoO8p5k+ej8M5iXJrojZDVZMzDUfEb+3wqgtdM7
EIvd/AMmG7cFdj5FZLc4zFcz02iAK286HHhmdkbyKhvMXbQX0GXDgiika2c+dfKu
kTt1xA5Zvo1EXPMTvYeSuBjgIWrhdJ8RZNnvX5CwQi8Iyzc8JTSBYi5tNtPXP1+A
RUphNo9SJ9hm/QHn9r6ZTh117JpQ6BkoXHsShNUBbqiDurIe9jJNlJZPYZ9hXAUa
Bb/8Ow+2RaNaehFx+5MBC0QvD5H6Qtsi7vbs2Yq/NzMT7PEz7fMUxVXdt7cvkkVy
zzKk4mk0KQ+YncpikAEHnzQCuP7t3FNVy+uZAXtPMGY542J0qSJK8s5IHpsm5wQI
v3d9gJP3kIL/prqL3oiKfHMImkj3TsrtxSs3cimSMvdyKPwKyrNmyeXBPe4sK2UK
sZz0aR8dUGPvHeNRwC47yutPC37wCwbjQTB4fdyHoB12O7Ai2Yvo6oybA7PJf9An
wVAdlEGgnEfTVDreQ/gYFqz9OE7YezD5xdg7o5fRLyeZeTB5FuecMmkETTnjP9xi
IfeGj6CFb19g+DbNTybWr5fgLnVMAqyMGWFasFDWy2Lo6C1iPL8KWCpejecMpf7D
vefI7SItHdHGW07euM29VgxEGs/h4pT2rs377Zr9L31ch39RsIjMvvyKpfxh87i1
ArWbKDVFLRKoj7IBWA0N/me4n2Od6NWW/rPGRSgupbmHpKqm0xSepyoFN/w26i00
iXmAzIC4QuyoTVOA8015mug3cGeZ0Rhi4+qVEZAyZiJHXzuVRR0yhsCeltQiLdWk
7qfIYs/nj1VFYyqHskQNJONUKZKmKodw5GCMHCYr4KVIwiF4dKqhjMx860c0BQx/
r1dnnyATwYnama3Ha//sW1yGqI20g/D1BpvcX60L1MEQje89xpAYdzrSqvuJfZZD
6gPBhmOZYyXDAZgxwYYcwsLM0/BCk81ar1u3FbR54xLSBTmTv1v9TKsxeA6wLXGV
SRQsieCJMUvZGsDyJT4tXvTp6sPea+Jvk2OOcueOwlbM+t+YMJWtVH9qwdewUI59
ZJ6d+duqCAPSwD4YoE+1x2HKdmR27FGeZ7C501FvbH9vh5LWnMybup55rUTrOVfN
KEw6T3MFyNe9G3IMDgNJ3AWR7dYH65AWDOu2+iBpbcBcr7uIHHzRS+rJlXrt2kF1
uXK/Nnt0IY14CKyy5MJqdVANprALn8v1QA1rIkO2KzILIAakNInHEUHdGNDV4rd0
sElhXGW99j7yuy+jvSyn20a5sxtxQF3Xd6lkfq4stwWZP+6b5m7gsgUZNhhHa+jW
cbg8YOO0F31dXWdN/Vy47dFC3ozT+eWXBJk73OKyRtosVd0ww+GOokfpXmIzgSQw
Hd9B/xPeZD6IMFfTJoy3WP8gxiCrbFs7ABz3BLP7MtHSbsgb7GGW/JXCHvbrq7YV
R8PWQvSKk+GaCkjSLMnxx2Wjd0XfdtDE1qc6zMQfO/L8EYJT/oKLKzEDfXgWbL4Z
fAFlBNrsKMX5/mN+ZEsbMgbbQmnwHAPRQUlHLKRFh0TZrXr8ZZylV1idmBWYDJbY
MdXHy95mgQqhVVUKgVDWT6nV7Pif4Q7pLLmHTOeE+HRH4sx5L7QkQ2FRvvyOVNga
B9C/663Vvm9UKLpjZBzVDY6FPRi9ugfWhLMxY1tpVpLOBDU81WAaH+uWCTVhg+p1
dfKDTbZlFodexOzgzrlOK9T1i0HObVim0CziCUNfj8eC95YF1hrgKMmI8ehmij5A
yqmZ00jvINEStsJul6GEaa80AXi5LGnY3UUz1IZOKApFgh4YSKZZD7cr5FCrHGRq
/maOyFefdtZRw8wM1QcleZ8fGDMZtRuNJGyFf8e6zyephfrcPRE53SnuNINbjpaj
bZMnzlHuwmQxny0yL8qbW7Mg8gdY+Yl6K4vdO1Po0fxd3taah/FxzFvFHnK74Mtr
yg1AT2O4y6C+HV/mEuhtly4mBkWALIWA6Y5aVxyMAavK/jXMuBSHFE2h0d/1wx8+
/glaRr4fYN2XSfarZ7GDEJqhDEkYmrSTYeaNjEDuGFxOzJAIBQZ/IyqRS82Rq3Nt
TtbtpRSd0mcplkye8HcFkriD6ulV2enGWHmTXpgxxuM6ErJujqwvJWHZGbzxoTR0
KjT3U/DuTdBrKWug3esSuzLrddBaAcuxN5BDpc0l2vV0oYqUonqJe1cXKVPSA0mu
gtXeO+khNlbiJQNGexpMV+nUGXP1x4Z7f0jpRG8bDgRnTqm3zVrfFNl6EZzv3xYA
ALuB3xiDkBv03sit7K0STF9eLCBWOGq0BXJqdcT74wZtRhisQRN8s3dF+GUr0Z3I
DunI7L+djPWMDoqPHMg/uQmRKWSCd2vaducTmlq9Q1z6FB7D4ZLtuiqYljr5BYd+
+phSzQuaw7N2/8Wqsth+6mhBaVWRC52grAZbe8Cp2PRIVl07jWF0gTLs9neH4b1X
hS6OS7kOgvxw35EDZisBSSvKBZKtPcSj8crZ2ethP1KPddgt+o/zgBuaBlUE6bOL
eQd+aKBeJgthHrq0QHSOSmGCCjNi+E7J9SWq5Q2DKbln8W+aSSSYZ4i4SOy60PKG
Lful+CTXSOyJTiwiyh2HpprYi5rreAzshNavjuNTZfCGObMVqrTe+6MeXDwca2L6
HL1+LbIKhV04BGJ1JSp+A4Sj5CCyL80xWYk7+1MJjxifOyIkyBliCCeD25PQq4nX
AsXIz0+VkVgZZTjUUCbeKYC9MCgnUHXOVbYyuliRiTgveZb6CrpUlabkVM97xE/5
qdZs2JKwpF3NjWN1zTPGWDg1fL4QP+8zjaUphCYCZtgWajWIN5UeM9kgIoRzLDws
JrD1P9k/lNUFWtvT+96GDIAXjJS65Zo9Z776FoGnFmXEV4xioIghOgpK6NAQJ9UG
JV31COv7o61+n7q109vP1ssnPCh0yUgW9DwZZkXYXfKV4Or5dDPNGtPGgf3qX7Bo
aqTlhWSWpogzeSd7Pq2UhfYxEpMjEthHPfOESwef5BgKiouZa08txIk7TyIF/xI4
jfs9WyHiHOaL/bUNFaEzdxkyrl7oEV2qtmtjP6NgEjyRxdlNFF9UtfymeH9E9hJ1
Fw0+vldJQwrIN3PEh2Wpr42EdrsrRUwcRHJY50F9n7uzPNHAZKeawyt6lCn9XGqr
CCLZXCDCm3H5dBg/OBndgQfzYLd1+6gnmEb9tU95cgHWHHWs+4Czd+z9MtGsYY9a
FVVdaKuFPQHgPyIOlyvRdeWAlJ/6ignCPg6WWEOLJkAkYs3IFMboOAQp1E/XOaUh
5PfPcF8ZB65nKC6ffJEiJKeihwRls916XKwjtALvo/oN4q94rssObgeu1KYnpzxO
nrP48UYdrOwcUPQjzoSw3h4SvQGtKXWY7/W4fXKtectYJvns85YQouIoRch70kRf
BNB9S1AZqIweP2CA7VjRZw5UmFhVkKzuMxD6wg3w6Rca/l0C/+Wd8kJzAl3mBzC/
AILI7beobg6fCNUdvdIbTBf8L/iOGveeMUnCGSNJ8oDdkJimLwnPbIC1OCW63l7j
vQxZYLpOq5k0qt0HK6QzbBj39q2AsdlGH5yl8Bs5T++52KLVYdhPg/8AP/+eyBv2
ErZ6Za5/xxQdwjM4JFgAJGgNZ12xCY0Ohq2CrllmJERWjzLu9iLplsXu5xqMlCn7
LyYujr+utLjSJoBTeEPQWUccPPdGxyeK3BqX04hyX5cSsz7aSHNItSOw3Q3Adbdv
GUaLtV+EP3dIQWSWQYI0tjFQKL+Et9DjN4doMc/S2Xvzd7/qoy56qBIsdB1/GQkS
Licv/vdeUAKKfgGSGrEZY2XPuDTXGO8pAg0a67TCo6BgYM/CTP4yB4YSNxsjrEA6
0E1cmaof2ARfQBnAPI3b2WEO9fuWs+vNKy70I+4eqUXxgTZR+KcIvHFKsOreAcIP
jWPer6XONNE5NBL2MZTkYxFMXmdcaVWYi6Y9HPa2WIQm1Nrfl92+xfOObO1OEtvu
HmayhhYpgWWA/N1R690Tlwziamlojfy6Efml36R1kzYSxwfhv7W5BGgPd/oFPw2Z
RT9B2PHc2eZJoLwRoveVXvkNVso9Pf31m+672K86KEfdUQcWhJIPtXqVyU6lhOuO
rjPJE7OMHSgGHsSJGbWQOamv2TuDFvqoEOYTfcyY2uCRW++v2KeSMtxuIzKpI9aJ
jNw8dy3N5LU/OYBfSYOR3i44Kx08sILWYPLW2hDMDgNKPebar3rPtWsFEK7yEKzH
doOVoMfduHY0gwPWvEeQaoZUeUWZp6qgMV3imvm375/KSlw+h/jU8bRPqZNdEnAS
Blnx0IIGWWKqRutCCF5ZGxbK1lvlnX50/eg8pzGBWcWnlp0OaPx0yJUI9UxC9Meu
lF/ocSLTVVsajwMu+jopEgECKL7FxBDDjgjgy5Cse3k8aROM6ekJycUkoInnAGuy
ZxaRnur8LKobkgq11VXN1HWrUz3oZmuPnDP2f+4TnQoZS+eIZKA7BP1+8NCYbA11
TbufaSc6ILRh++GmN2jWpDWev1e83eT51pyOMYl65YtFXk4jltNZenF24RiIKFYi
Wye2BFaj/rNhnn4PxBqqPEzZOroDJYUDcnwJSWTfvkfi7nm12kRvIgh8S9BF7Pb6
FEbmJwv9BahEZ3Vpxzvat2k2hf1zvGwyAyK163FE/jZVkO2PA28tBm6hMuDF+u9S
DwapADKSwVpfTrBm2dYgsl3+nyakDr6r7gvwxRcqVv+B65e5RUJ3yiLdxxYNnMLF
Qc7bveEbUKWelVe4dA7fzG+2+Pl26xRcKxDEf71ddelvljO3OOzR+mAMFLNTlzae
j/L9ci454rbONG87wgbZTy76esVtLrkMBx3+hUhgitEYWd8rYU9YCMUTZ1c3Y3db
y2hYotTJsF+EjXMEU2RWBxj6IJ20RvMLS8KJsmu1GyGETENf5K8CgQW9Ao6kAsev
jS1IzINIuG7gC4U293ZI32omo5mWkY2RHE0GyRNHX2jnopA9R1JSPo4FDQJErdBC
iK54R5GR1a7tfKvLt2KiQ52764TkX7S42Y5PvrVxXw0UWGZaf6FHl6YdVGtZZH3e
7eEo4T5vkA2kWny6RQy73OfRJ0vDa5XQObpCcWLd/aPI8yiD/gmqplbCJ8E9xnQg
amAtw0aAaz36jcBud/p5jLIPIWu3u6+FJS+qyTNsReEEwvIBJKSTtCKBkBDPVUoB
NKUkbmxS3BiRAEp8rJTwkXZyxybAPnSJtlmSMn1i9IN1+K5sTMpwoisGvm8fC/9W
SrtdBI0hs+alS401xAmPqb4+eDHGK7N7fElcrcISMOiVWRb/zwI2wc1vDoSKjyM5
0R0qfloEU6BEc/Ld0FZqFBv314h2efi9rTxRn7xpWHqaUQ0qiJwTixsJk5RVONqf
BFOIZPX57dFJEbLwCNwZQOe63Y9hOg6KjfKmENIfC4BFRcqpdyhXk5JZ4gMOpuwS
PnK0h3PWOFzwsFumShgiXLHTbAogHMXWnIrsgJljzfgKSE//3SkXCj1HcT0I33lD
8PeWIGb5pG+lpP+UNKXCyw03OUs+KhIY/Jbd5pdsldYOA1RhUB9RQYwn3cx4rOGW
kdQVekfN9WWfv95lRnUh9nYWqrSFnhmvkERARHVPNQfy423fsxVSDUmfrmfAQwvA
mbhmFgTGnG0bYxCMDdtqeiB4b6fK3Yc3wHcSdZtGEvbTIW8ZLs2+YWdH6RHGVDRl
MAhhbQWv+MiDzL/IWojwSJBjibCQtxSMhn6Sr/GAN0B8ePbnyEZ89Ls9OwA1rXas
dFOBymyFPi1pYAr6sUfYW44+n818q0rY6bgnkG76vJXc4GIV5yBzxcBWAcQk0MUr
UWQGsK0sWC0orgUAurvCF1vWO6JnnzJhI6qnE4KrUjsyc5NwRUj4rqZDc2Jw7Yrg
mvHWXWWxP+t5N0oGcEQOFD2kQghwjV0dbgy8f7KrjBUqZCHzX2zGmGABTgXXxG1H
yct4yMjYZ0CjgCgLXZBgGvcPa7XaZrDa+hH4NoB1rkTZbDwbc1V/46qKqFsAjWRG
RjOlPJtun5agfoSQYVFv9Ul90Lx4iH3uUmk8Lbt7S/HFQziz8qbfgGn2asJCCNEF
OXUnFSQtffd/w+m6nwAjjevkHO1VTWRqVTNLIK7z/V43oz9iJNOMRDjZA/se9KWU
zWu4Hel1+sAsLhQzdrxDI8CB8wHGCfsilmXxtpAhYz7GKO9yf1TDqhgAqLzJksK8
gg3Dfd7CBIfoisia2D6CAKHKWUNRiVokSy0RCD3SnZAUiwnHhUuNZHIwaN3uNpDp
E8ap6U2CEC4de1kuT3gpmKi+LD596Zn3VS6IhGaHaEp8zSsHcT9S3cF/NVNHaiV6
MFyRGjSRELGE+R96l44Iud9G7iEeyd9cycI5iAvf7xNbijibFh8uXbPbKR0cnzsZ
9hhSJHU+sk5EHM+l/OKSeHFOHx3GqC3lYcFo20a+Y7471m5b+W+544pJlURhQdYb
h43UNddNlvz1HlOHNcZ4NloRX3k5yuFQP2Pwkj2NvBl+nPi2kJk2RX2rnMzB7OCE
1BSb3WClrZHqpPx7EiuNDw8pl/WxPFtoyANzkGJC5j1f0xlhKvFM750RMVt8YzBR
KQ2IFAS/rBR+RrD5LX3C0yrmtFx+Z5nkwa8mwWQywBo2Ai8iAQX9eZHg2MXhs956
z+42rx/ceQ0sDJijBYLMuEfNiEaEEUpFpdwSxC/rGGa0IP9HcCsf5R1vQG4CWcAM
T4UQBJnw7KSbWYeZMZLwdhmMkZUrWwq9VPLjXDf1V2ItXzDnxXiLSgSAFpmj0AHJ
dW/CPZFokMYpXjbcaCxSW2fgw0llLxGaUoww8U7X0oneBfjLGIngI9k6zXZxYIbJ
nCrMwmaqeQdb7S6cpggGv0MJNWE3oQlhBTsyOtRd8/WC/eL8bXereqV74OdsUfpC
rkedRChlwjX27BHntRA9y8O7Z7GTVZDibT1fHofKrzPjoHoKF5/DRc7T5Z6l5yJb
Vo6kSrjy60XZZmGNzcP5rdSiSeFpGbqgs7sknBgDp3houCT7zztuGFUAfN1a65j8
F511uWnDaf1qnStkeUG0fHQjAWuQ+zkluw8wa1W4Pn7FOdpNuknLijtUqDbGic0r
gg8nkecF3fUdSNIRKVJAC9O5qnsw6rmMGTAcFZx5oXxCabeSriFECPdyHEX23+mK
ghn3zncL0hY+CYcJvBBaJq492T6q6ec1HhWmHov7zUhDz4LOv/Zu50BVmPqVsXmM
Xt2lwSimJOXhh5zAA7/TCQthFFru7nPtG3bVLTLdzoXvxH9WJXf/vhdM7hEC2lxv
LQPMxHxGfMBMpefodeK94eq2+c5REgd6Y5ZWE41HoqUns2wgoktE11sTlD8iBME3
gFLgBkuwGAChNJMyzgfEtB8TLrYW68tPbuxYUSMRfRMnyHHjNaFsyoa4QADVgTYT
GqZ2Mx8TBr5G0VePR9hhTdRy3Urt3y5oqyoVQGOPPAwdfHCkvVNqjLE0mup0jsTI
8/6fyPDaEa1J3/M8OFEd3Q6nNP+cl7Vz2syJ9GBmct55Z4qji5nMp4OLKB+2mTM4
Xx9kfLn3fxxBpo13jfgUOQ9AGTFPD3UeJS2BbPyf/wUajRm96F6rbAX30hVj/FKk
Ug20/li+ygie9JfURPIz59gdvHjYZX4AW+Y75R31+mSyeC27lTmbj0McAD5RC+33
X8pLc9zNmBf1Rr5oJOyGtTB5Gvkt6k7hf8gnvzr74GH4jXZV7c35VGDWQ41EJVDs
4tSBeKyRr3DUuxc+PlQGftF6Jogt7QRYhe+4NmSmMXwld5PHoatZhwGIZf82yuoq
JzUcTIePLk6h1XQcG1kHEgpxlAHZZvj/GvfEAvY0lZxuVa1kwmGL4pVAlR5i420A
uDMOhC56Vy5P8xSoyTfhfqjDsygvTJxGL9nQla1xwMPAYNvnpPbtMTSlGyVnK8Ib
UFXk9zVLY6J7JGAlQY6spMe1Z78Zydw1jGhaq7mWkgVWEjZ22EIu8CUDN547yw82
ZM6SgoD2FZSRwrwRFdBFUrbqBsTPQhXQMxYAMR+3PUBPyEClgoFKpB+ngXnVC/NV
64yfSoDFETkbLvlEXUtWTNUI4NBKrMX/zpH1xmGc09doFtpo3MFTAsMkQr1birlK
A5wQK2pZ6P+dajFFowksppTpbZcn4sIDzAW095kyhIFfWpPx7FLMhylpnBt6e3Pz
1tSJ5Z0ijTuU27b2cgY0gcBAzEz+9MKWKToUntsZGUPL/x6BCaEheTh4pkv4/nG0
kSk3b4yW881QQeqUeSPG4wQOAqdZD7+AEnBAA2wma2glzhzx5Uu+x8XyfW8nBomA
secFLF/t72z7aCBJ6fzGjsjFLEL69xIYPcljZQUQk2y9YI9mERRusC4vN3x5XHyc
xpiYLYFHdsIf8iy+tuahMccH+I5gjkkm00yaQhXmCTn99zfpc8KkAm19q0QYiV/p
LdXVpSNtBFLcJDEy2T/I181H838f2gj8z69enMMnwsFKYqvq6UwKgCU6Lsajzoui
a+TW8eOmL18Ok+vT8uoy0AMzsKEo60Ez8aqMBk+bjjoUiQ+mgkZlFwIxvefscOTD
oBYN7NHR5bcY3iblWL5P2CaGHnw60aMlFg4D+zoCHdpEGNNW89cXGSB9Kwyeku/C
UU+IMEymodWxXu0pwKlijRR3SHZ5CGHdM/DXkKmLzy7Qt8QOoRhgQe0CVmLSgsGL
JHBPzOjIDm9KNu8LbcORkszUes9lR9qX7bZYPONreuYIPFQ5Ad6kP2fiuRptLTl2
wClW8QCxvQRM0TA+wlLTT+kgUcKsyjNYjQj3RehMwNMGcuaVuq1QuLW+NMvpO+ke
7tlLglr7GwtqlOM2MxD4KpjoV1KRhE9qDMsAFatKNHfURzMUC/mK6j4smFaRJjcZ
ds9bSSnUrr3Lfw53yHmM6ZXWBFh2tyObopTQjNoMpqvjWH9lIkYCNBUHigdTLrw+
qDmc7ItqxPzuX8F4AX0+DQAehmp6yRSiBzNZVaKvXJgGsCuWBC7MxUkuM2SgYEC9
jMv/uiIlFY8iykrOtxxhgHw/MWKEBw3/802GB6tY7fTvB+cAoz/2V+zhktp7VzCG
b4OFnDqHArpKLUa9BdsgDf43L6gfRs4X1t/qJ1nWI7lGDQR5GLnv/agrSJzfXXyN
nt+hJTUjdIMGbWmc/DUDLZm5CUeIDy/FZU+nLH1lOXHKbRDm7KdhdIcpDgPm+Uwh
RWfVDmS7cY20NSj/MhcA0fc1aEODmh25T5pd0qmMOc4me6P/3Ux06sgGlCU4UQKQ
ID2beeIk3frVslP+YC0sgqX/d2Y8ovo2OngzDVz793jRj+/HrBA34O7TvEd9lKdJ
cRQDbxpN/+hzk33651QdIE/ucwSvJb4h46SSZi1ZwlCbTr9EOAwvdGGZrkuFm8Ko
3XHwDiQqa8o6eobwJJRVv1Qegnwd3LjXOBqxN4KW0CbWTtQhVwj3NBWuEbGRtDji
elnyn7Flo0sspfFN01s25hX3dAwEKuC34/YpiECGVAPMxqptlp3iE6oNlShlBmA6
ya2xKEpg17kcmQA0Gt9wgpFQtAIQqmsdaok9ylqAF/0g1IWHdMCEXcNe90fcgrU2
/qVEOAuKvxZj6sWX/fYxu7CgGRO7fBbeR0xUADtzfEYdQNPPI+GedxYEpNKiJ8GE
yBrxubrASoNeXzJtvqerVuHJGP5r7fy9LH3IeOreRObotMT45VM4A9oOZSZFZFIE
OgsLMoUzcssc3f8uce1fYB3Ntb5WuyNrGVPVWfUVhQV9nkUiF6silj2XxbGUH1l9
S6NG8oJoxTBcGOxPn0ljIjFHQ4WG7t+nIa+THhBxqqVHb4Zoe7c5Uhq0Jxl/efQO
ucCZiHbKEOMOFkT0ZwpEW74U+0EPDpmUXJu2l6WoTmV/kTQHKK8nLMD8GpPAMW0c
JzemOrURtN7hbh2jTFx45o4rsZiIdY6Ie0ZUGbSqjYghPxzgXRgRa5kI27NNSCOu
/TmnOduHMCQGP1ggHhMFqekeomi5XGn9073IR32+yjPR14OBjQTEUdXiC9FQmGTn
j22mJ1QwIOPAqKIwwcT7mgjtXZhczcmhXowtS4CP5Ghs12n+iILnQTJ4ITHkqmOv
iQbsj2kJXJOK2wMdK5+4SEliQDo0YLq4+SenIEdflmh7uwVrtIsAk32O766XOVTg
H3LmsUtOzrDKQB3E7VZBo1mQabrIgdOmON1CNO+E53PeokVuKudanh8twxIUEbOB
I0dND5MCQiBi0lhNnBjqBSNqQbNkexVCYhRx6HYd48/wsYmOCOORVDkIafVQZAoC
gl3BXTArV+qERXZ/iKajTlGeIoZ+UxDdZ+hRATrQFcffAwh9oXmgGeDhC3I3w/yi
HDukL5rOS/PYnVJpTceL29tjJ32UY4sCLgZvVCW9mNSIB6PZ2FXhEfIcFpy3Itai
TBUx4Fc66o3ag7HLccEi0R8wjMY0m8ev7ZUt64EWJj9EgadkrI7BbHUD1afjw6fa
HxTRp2lTi3TAiGlUpBPK5ILKZ3d4VCQ5niSY20S7BdIBwDNMq3zMci5N2VvZ9ypU
A0w3F+p2MBMx1PbbKuFQZ8SSYPcLgikccaftT7o44bXVDd/jYcEs9VQhV7ytw93J
ILuhkZL8zxAgjVyr/3Gq+QuDuvCe++DLz7bWeqmC6m6llWhOuLBlCvs+a6cpamyr
uvdwZkq6xo3sfBvbZoU9l/+2UJp+BIlKOjpXc3Gwn8fPzHEYdnQ8V7bNitZTPepR
yaai+xX+0Pi7aVONUrx6OFeMnGOiwLl51w477UtYTFSBGAo5D94KycRUDDpiNUMM
y/Gied1GnYYDqeWt3tSd39Zl01r6owaXBnTtMiEm8xnz9v6YIBedzkryofVE1ReK
M85ljVpnSpLe41XG9NZA57uCxSo6aekq8ZE5P3Oht41nu2ZxJMO6XJ3b7FMFHYeR
LEONpFXzb2wwYwbdZigSVsi6jvTKAvrQB8lNIf1YP2FnOBwBSspDJRHEobTI1Iri
BUW9ALqWOjZ1SU86DmmgP86lyT6t1q8mn3CJN1tyNzY4Zb/28LxpdJl8Z4B7NmPV
yY2O0L/oDljbPYPM7nPGlZ3ZhGx6LBZysvefIZIkn/fya0VhS3iCbZc3P3uDY9xm
UnSl9a8vEhbnYa+gQfAAUuOU2/VAkScgIp1tz85DxA/ylBqE7PnmXqqEoxg7f3K+
hFjaTykzRxCAT4ufbH698yUzVxnIaTbWAPjFZl4Z7S5m04BZNBbtXAaipsoEI/qS
QqQykLC1Sha3OyKXwvg5He9HgF7gKT6D9CqyDtyG50n+7M9LI7PfZYn9GFkObCMk
bwG6kOnEfClTyUs4HvrrkorLG/FpWkeXDwV6D0wVpnYf0gbiamaHLZz8fzynP4J1
lg53gRLv1vxT+lyjf0OIVqwbncCFg4swE534vQUGpgB4+n7U0qVfN8XjSElzpEjA
3NqQMSUtkQgdFHnJMuYH71e0TpLEbeH3gH58KABy+QIziA9eML63Q6p3g6K+MzJT
c9z2e6kdXrAaRLKpRKDfoZWdLASFR9be/JMczwWiKIUnYHcJ6veoAH4LlzUTjpFc
+xBfU6e9mOXcJ338iiSIqH5/+3VjHmXtTk8W4TF6hHoy86XG2bWU0QVQfa/UKGII
mGQ03VE1JAcuqaIEx97LVlCuD8d2iuX0UDrONjn1730x5Sxx8Q4Pw6khyg5dnOtr
C38LUS+0hcU4pQxadT1RTtIURPi8ATmPxu9JqOfFUEzvswN9RHKlOsCcJJnYIo98
qOJG5iISSJuZ4ouNhhebYwwRhX2Q6oaYSM++I5zc5ISlkjFnAX4UMT+NlNcByGXh
9QjHz3jlJXZGsVxXbeqnGfFMrCbHq219HUw0d5E7JrA3FyBUYrXkQcHldJrEoEPV
550xiBR30CHjsGLMJlHxakTgZDswVahWZHk0Jjw5aPEnCqZCUtjMfsFrSwF3AWfw
DgsdHQGGxM8dX9MhdjwLp01u+Zfieo1Fz0RJAzcndeTHBmKSuLQEtZWlzJMTpY9r
t8deaPFzAkEyrhg5XhE6O1kQljMhlOhy36EspWxikL736vRyA1BpYpsfRDAUHgQY
W77dFHrVkIu7qN30jnovjq74U91k0wYvbieDpzwJMXsi7AFJlKrESuLahW9OUQUE
Vw7IkrDP88RscXQzOpsW3oyD5rUiZc9ut6PzuF0tAbsZDlEmhkd+al0JA4H8YCg/
UcvGa8K+MjKmm0SM/prgYQ5PL802xsPeQ7vT4XbxCLU0fSXV1kfb8hkwaGd5+faY
tUifMx7NtqG+iuki0gqWTTtKTZV6/DcJ96KC0t/YP5JGuElGwP90lrwiWCy9vizB
Vpjwcyshq/avF2YOTH42k2uAV4cyDjiYEKFeb+O/cqJgGJBq76lbnDrxUSm5n4Ov
OtJSTLFGOzutkyO3uR8p/BFNdg8Er594MA72fLm1ynVWQzrvE4zy8QF+CsO6n2C9
1vibRjGRd8wC76nLhbgES2R6xU+oM9hpP8hU1k0SJYuYqUvOvfx3FOhzXLfOddlX
B1iIiQc/kswVVH+J+BQuRDFMrximB2YiNzo1ltQ8z4+qgVqOoUEPA05rAEiBZ9AO
EV8kftmvIgHpZARCEhNChGQ0RU2a2b2PQoqb4krllzMpuXSE4ydcMq8etU5lOBwe
52HqNigO1f3pvDnqqDRoOB++bvqtt5AVDvPmHUCWRNkCAnDSg9Z4AfP4osm5mJ8h
J/WLppXmh7JzUR0CMj2y/MaPZIELbkQu63hXkJDDMHS8uLiCZ9QXUxak+uHEThwl
GvE1sSS9D2AuKjnq20RTkbqN2y3PVeq7kQMkgMHKJz2k6t20Wkde5a+grFf3XM/6
0fWVVPtXp9xhQJT3jhB7hNVBwJJ3fPRDvROSW56JoSPmSUOB7OMZek0aaWxth4+m
Vrf5gVCpGsTmglOP4lJiN05TD3Pdn251Lxxkot8vBWOYstcUWvaa54YFs6NhEL3z
HPNyl+UZxxG4olFb3RgaCdkz35dX3/madl6kKlHu+kd+JepD7n1bYEByiueiiPf1
hh6oOxWsAREoJRWlyepo+vzNF0JjiZVzhvJc+1wCmRzlcdrHjDhDK5pzHC4cmZP5
HyuIuIjAqHviARwkCFNkjuN3dz1eWNM4FNjrc20YjbG12i08v/T6j8KG5LymWuQm
U4PnIATd+kRtrO61iYr26DTCj2+f2EKu8wq2+MLBPpsR6/YcSNjZvUG9c5/wdbPA
KAyF+NSe4zPB98BaFK+tUpaHTpQ41W/ZQkBhqdrUcg75B9GrXB9vTu+9pFxwbg4v
OJDlOBHo/yx+pM6khnSeW3Xh82z+QIH4lFQ58C/mj8z/LEwUoxfpfUJ8IzFT8AWK
hKNLuUreAeT1ajPhSjm7aHaJQgzuDyZ8tUSuoVFTRSqxP170WddNjQ5P2AR7b2PE
XX0+HwGghUBYIgZW5Wtmb2rbmhj5VsHIe48z6dnsF59ONk+43VeDY6woYoaw2drG
1CnHPrMMV9P0HvrRal5eBSmHbU73E0e0wrfzV0UuYv/npZi6n7/tX4A4liatyqhS
gSAK5SGUSowGuLZDVgxYNvf4oqo9RndmnqAsRHWpDo6b0w1VMS7FtJwP4brWVZbu
sN8nkOB+8IaUGldcKY4BeQYEV/7fa9B6Nb+XU/urErhmxzU485Eb1SMMDKnoS25A
CxSUwuUmrPaCI8yu+q8Yh9Hj2L79MFVfK5Qhs3yu/n5q74dzH/KrV5iTbrIe0zUD
zPkSNRqEk/jv4sN1TULH2ObDxk1z+nNYn4GmWrDLUqoEazP/TdaWy2FWp6kGigQx
2Ae6/iiLAieGtmDhM1QUrQazLv4KOimWV7sGTmJVVYeIDuDjAAUy4I92dXGbCdGA
xKyWJKGvtOiRhfkXplYgWgwgzONJwcMzwolR6MhfAbPAigsx8xTicvBb+fg9tiBr
++w+DHQmTVyG1W8sXzqXqRjFaJd4Wnp7nviCkm3Q/bG9duK0pvspKc1Ha5hzkZyr
uXx6atraEzK22WBIGZLDppKSVTn88xh1FnpC3qioZynXAcyloMc4o08kstoBiyDy
MDTSbVH2tvSUg8t+H+81Et2kS+j1xcegFhg+y+M3eM/erQW9axAZxJuarzGAHxAN
8PODAAha+jDSERro3dCZzE4JjdZDZ7YLE8RMVOpBE+NehrSE9Hs1NTvlQeCuVRRZ
r6MWiC3ZSB1BXEtHxHxfyxK0R9h3lXYtFovfz6qL3FuX+2G9rSIHXDqxo3XeRtXP
MU+Ci/7BBVMEgGAcXl+IaMAw96o+IodK5YGAqR5rs1ekDteunKhf8gAq+9yQXxNO
x5zIHYVZoNeexLP89O4JoIC7X5oBqZdBSYP6KytwANE5YpT2LAx3lJh3LmZNHM7W
MRz4Q7PlZqoVHnLNOSibVqEg3HGnUZbZR6PHvLwAvoYy6XBY5hHIrXacaYgGRvFo
RnWOvO8dxKX5a5qgkJVl/4r8mz1l8JOzShuS1GkEjFSswPK6KLMF55oDnWsp7NDA
20Iu8Q6HVBI6telkyC0dyWJd9f31TTTsNcWmv2N7RyejjjlA8mj9jVnNZReZuM7X
6YMEi7iesuwV9kcKbK/y5+PaO27mNJtVnVkGQ8KvCo25hvg8ebotkAwS9gvHS2zR
pgO1AZwwjB3OpFPdaWzqjDWtcmgGQT0k0IBWcG7yhcfQlOH/IjwzFV1z9E/1DM6X
sOz/5Bwu/CNGyxCXSpcwMZjr4Dc4iC3PyTpIQz3NLopZAZAva7wT335VliMWUAd3
9DrNgjL/Dh5lZZsOU1FvwIFWogvfzye71xSQLXyxlc2RSb0iCtWf9JD/4b3Bo+6Q
y6xo6YVH944BXm+c/j4ca75X08UIwxSMybqiy7mTbGCN2s012tduYAVw+7QPOpCE
XvaEfLwP4S8+0QLabT1UMFTDxp4UujG9Ob5/9SYTH9U1RK2pdRp7J4g8Hko3CMyQ
mHSQFhqS76MX1ZW7qn7NOdFVMe2Q2qLxPNAZaBakgFvqsC3Yakd7zzRlw29EB9OO
wUgML+9BFuR/ZUUe0U/3cj2oz7OLzWO2xQ8nSDxhgYn1pB8kjRgRb0iEGkMy+oJ9
4tQi0rqR/l2G3drRnXrzqbgaCzxIdb61G3F2MBTIxnhbUcB0XL+jjP9kQJOT7xVq
+uPgZgpxWqeSoTxayTd8bTqSSQGkeYa54niASF1JCfF7B46fFa9VzgC+/lN45gFK
1d491j5qPiJKNBeeS84/UEqAMrM4IHdXz6Y38evjbs59aAwVMj1+N/0YUegbDD9E
xQNDxT5f91D4LU6lQw5Lr8xt2sPT8wdt8fHRLh0uLCeh0GQ/W31lKxPY7eaeoagT
eZGMOdWa3DhYTmL+MCxD4anYlNi58P7Y1aR0Uk5PBuPY1Y3t2sX1YX7d/mZX/Jk2
+7bGJKyt0i6NFMYNZ1ksHvgo40UlVECu7CIHvBQwUsK4FAyITvE6SehaWs0TBylP
ysmNI7lAxFqj28b0MtY/1Qs4Q06U5F5+NK9BqAViM6EBj2A37p4Wjc0xrsWVru2J
iL93OTAQBX1HwZpweQzMuenx4dXmiQtgD9mNFNna3ukv++mSmxdpPRgbssdZmY8t
HX6jdJ8S6hJtQv3wRTbKCnlEUdiJfTzaNuz+wp8JsaYxFQSg1PRS6PrjGmfo4LQX
qLAM+5M9pIJKD71LuLeZW8ctsy7MpXq56Kid5bGukxeMWtr62vxt5WOq6Y8ccE2i
BfmXXWd6HEgLKPFg0ZgB9k4yKs8OCgR0GVgxZdqlZfw7mcViGU3on3ddW1Aq31EW
7WLfQsH4vTGWmLaH7lSWPJTBZIkumGfFCp4HgW/VZo406wgzYDAioa7p+PtxXodM
xvLyB3rtg5zQQIVbdqO56ZC2B1YVnj8THaQZ9A1hmJeyPpQ71VHSdvEzqzxNyIbz
u96G5Et9YsTmkitJTZqYok+cCKCwKcPHMIUfT57UPT9uMHIh/XNE0rOLGhpZArxI
Ekjz1DhklIzu0KcAAbox9MqSbpYOJI5vyHsfhj1lzIzGH3VF3/HmCXOW6lCwGXyw
eJzvsrT838UEqwot3z879j037Nu8ciHXIL3xN8CMSzm+vPq1uSR8uk1wh48bIQ/j
AX71gBHvNpreXkiz0Fj3ELzT/mLCpFA6yP3cSLN2uJmqqqobOryPvT4nMbS5vEii
AQ2SlHnWsbOHjer5Qo28ep6nIQ+tnHUFLpkVUFum9DXtK9xHRmECvGudjn7NX4Nr
qfNiUdcWOA1sJm2rINssfUhVyWQUE7tjAYLWeUpvk/KefQk43f5CN00V8ss4TzvL
jUQf21AqZhaf+EbR0QLLrGToUPsGmZrdhfpaWfNlw9u7GP8MP6RTz2xTX7V3sHqB
W7riD4emFXhdcawgBQn84ejTQE9o8Nf7vt3tx+FdRaMV/8b4Eynv0s3XKMPHeaxH
gESa/assrdXhhVp4OoS2RnosaFv8WvqvlANIGpV2FmhDCLaCeVdG6mK+WPHu7dGo
9t+wxwWojY31+DjU6/9k/pMvhc7odMv9ZI/w6h0buD2ucrCj9+Db4E1BPifrcr38
JU8jeWIG13/8Y/J2P3lelr4iP7Z9JP05uVGvsl4djxhtkBqexRJ1nebsxdEI1gwZ
hOhdrByHBQm+UfoQwF1uFbh/V5D71fKV2JhtRs8gznv5jngFrut+sLQQjpiqLr8F
Cr64bAhDrB2m2pICn46fO3P3CKg2yldL/mA0CwchKgMUdZgvBzdZub6zaUJAEv61
+vFBIaIsgGGQk8ALshSvjR+mSEb6EGptcHSF5eJs7OCu+1s0qmutXMFuXJAN2qq9
2I+o6/MZJ7iHCORrfiavAt/AmR9Y4J+o7a+cdceEgj058xk2L/4B5e9xxCvzq/5j
GBOaMpohtcH8mccgzzMz86JEqsQLGZ7+4N6TvPPCOeGSk52n+y8Mq6mu2Q9v9t+8
NF0Xa7Ty05HcqkWMZzwo6apTdpsa6uOvi7QYvsx9i+lCEqk5FThEyN7hKSakgWuC
TdUzIwBLtiLNY9gCtx+p/uOP5CbTkOjuumYZ3LM/VF3PwQGku3ri2QYIUrXwHVeP
XhFehTobwthGB23R+aEgTYANpmpFXhMMqthDy7bt/1aeAchgYPsdz9FMEP9IyqiV
uoRvF0Uv3Wkateo/0lnav8C7CNjUzA/9Sx8HyP9+cZzIqjPkpbIokPZ07lFCsWFX
nEaRBavzUht8QGPHN/oOBD2VY+QjoXhd0qBIIQZb1M0vnHYA6IdCu8xDLNzD9s5x
MDApau7b9qiMBw0Se6RO8fooxj0RVgGZb4Kh1SnZWdIPxtKvDV2Oo7OGFi7iwQze
1wvlvDfRrqG2PdYBT0ipRx+tjSfb3AS9D+cm2qu+E7TXRLA+erHSlS1sPzdGXIVC
4wUO1eL6vuCIAPNYfXHWxkpXCMvlke3YgrWjN9vdEZAuze7n+CaC/D4ep9WXWWJa
FKgngpTiu29rLRjGmHQwo7nGnzGHZL69cNZT3RokDBfyc67FYF5NxxjmNbKFaYtn
uT9A5EsY/EJCTSHxHjNB/2pDHT/KweJ62v7NC+M5c95m5GdEZeCkycLk4vhm2VrQ
KNbEKSD4f1D7Z1Ea2pim/JlSZULRure5k+OD+wQrOF5P/S/Z4alhK3fQ7p+zjklh
FHbDWGSetFbth5xtRlaA0v2BKRlIO03RWgO1ViynSmPYBL7UJMlktbYcL53N2Dp0
lH72wVJid7jVJW9m5hB72EA6t+9Ex8ov9+r8OoMekeYPhR98SlOfHnXiaj3lVVf+
iK1DAAs7M5cRVJwQML1pofbPeIWV3fs8NsldeldVo69/XjIv/5Q2xiXijJ1h2YQB
VV08yntEkJMj8kdB9H0peI7yskHUcDWtNlZiKVr4Uhmi/wUmmwNuuyI5Ck9smpmn
QcagsR55Y84YgImJCejyy+qLGTk3mtj2DZGTFWRFAbHvcCDsWmQUFDeW3neK9nOR
D3NBYi+1CYYKDRWKcrse/ugKdNfw5i/FK67sd9CG3pXnhA+d0AMbHJybwTDiSafI
V5S2fLYuihRSyzJxUgN1so2E5/TsO4sty/2WXIJn+6KK4+fnADz+CAoRYEb9D0Zd
CJiDBLYaX8H5ur2eg0MVw5K7tuDE6vr62ECNiGzz6AjdKA4whP5jVLD1yrFZAeSG
8OpfUVxztccb9y4VoGS3eCaLkqObGyfHUkkE6fpbFsjBySaCGOrNurgC63+uwJal
lfhG9SQRKMtmTErfvldKB6qNGxP8V2CqqQSJ4J+UGl711+X8togI4LESEb8EFqFt
C2/P2+Q4ou4jtYM4eP4aof15f9gIHDldaQYyXnB9Q7p5YA8fp897+pVt6qPxwSJt
uYCOmcpTfd0kyCVo6A2/+2EZigy/96uYoFIcVAYObMqEPqs0XtpghnNTwVOXwDui
AeEMoOA5uUPBsqmzcnS5U+HyuSG/Nw7TWOrb6ApLeOFmsFn6Lpn9U8oppJfBB4M0
xTvzBZVdL265Qd6Qj5+gw404QoC12fWx2ppbDjtJcpAq3Xv8G4GxOMzyYu3Ud6Zp
QEByTuTC7OaHd6c1pK4fAFRXnqjXTVUJy87KSEwC8hCnDrN6ZFweyL1A6q98z4YM
Ss9m39HR80KFsr7yMvFQTdCRrRChRIbcLhkoVIcy/n2kKdw6Zp1jYRT+ZgT+lGwi
tujlZ1UhDZ97PQgTt/lcZvW2vZVBmgO5UmW8kaoh0ZHwAGwKj7QIRIzANz17dlrO
02M/rZ2A4/BoMwy88y6VxSkHQSeZKKV+CbYsw03JAI64MaYrVqAQc2muBbNulXYy
q6Gh/whzlVined7+evTtZOlEKxIA/v9H9k677cFJdg/LF35n9kvtKgvAm7DCKLdV
rk4J7kEp6uAvW+RWBAj6yh+NvMuA/8hXl55HBv3V0WyqywnLZRT7lo7XEgf8zj7E
getn+y3bKMEG6JJrrGcCT/ImvPu7W7/y6F/6P+CN6p/fDNuV7Uty6qSseP0fKh6M
cvegGHzAq1hnTMxrf+uCz4K12NUk/lurMAVUq4Eok2AmMOxdTvtdFaUbWWWIvcHZ
z/QckkqZUOY+5CBUHEUnPNPNR22F6bX0+eWBmw9POmC1YrJkJYg0p/RhK+jPllgi
gBgCZs73af9Udf0Lv9vJi400RirHK/zQKgCIB0gC3XbzWP8PQ9uugMQzXxZa5N+O
ESW+wWHdbEu/qoJpO8169vtghinDPcP752cUNtnlzmvBKjTup3Ep4rY1TE4vDBan
+8bUthZqM6C3k5hAZy2RQayihhkkVyYKkSJmAxStv8rfMm7wkq7K5qeCxXGqNsCB
AUj0dkDaJAXHMBzpJynzMwRLDOrX2WMOWNHYm9U8EEgBL2tW2c6TeI/wh6BbtD//
ZZnXBbDtq/hvkgxPld6savdtPs/ZMzfHogrVIz4yqpY0zfA7ONoofgFIsn1Pwk9e
LXKNKury4cyfH2WSHfKVPS7f7JCgkENfkJx0zAq6O+YZIVg8+azKPQhdvyBFnhA0
fuOw53GlZaRrZKktz+UuMze6F1roTGjPe7nLSlYjvs8fBSmv75OXKxnmuv/qr15t
QK/9VfHYyAiLS92TJzV30FEHdQFJzHkeIf5XU76fQjIXpCAWuB0Ftfo5N7nVEwNx
KEIb4l1g9u0+LCTpuNZeM+G9RBDe3eDFr74v2bPhdVjlE8f7a1/Mh4u94338E+ZS
B28pSwK4WGpiC9jmCVQej92at0OwGTRKgozwTtAfbAO2V1Zu3J24M4f3lifd6NKI
EEL0YVd1mGXrOgHv/LSw11Ch5qWUUV7iHMZsM9auEF7gTXSB5ry+X/tntXiAuIcu
etyTu6Xh08jF+Xic5TUbELCfzH97KWwlw+zr5VZx4oYHWo+nmHnV+jedFvqo7QcR
bs2uZoOKVUSaOUuWR1T7J4hIm2CoBQRqU2bTf1LRn7MFgqXGkqFS9maeuWAg0Q3S
XUQgfdScesoa2rLgtUSR7RGwm5lumlTD60OfTMWYS8AM9F1kkNNsGIzxI8bVlxZE
FWtyFHzv47MGU2UGYnbiSGE2N6+3QV/Fn6M41Z/QFZ9IFmjnApKk2ltP5/IU9qZc
uWg2w+JvcA0FLBls5aFQyozhoD5mMoIRiWXu88cv1P+A0GjXMlQ82YVz+ajEu4+m
ri+JKVJS7ZuhMl6gyY3YysRWPcGdL4QIBpO4nkJz1HztT7LzMucupT8TUvdjCv6H
+Wg1aBCuTrpgtoe+K9XCxKQz8nClFPkN/Y2BN1Xl2mpXdUV15SLUA8kInQVg3zSX
nClFSEdbOSx+A6oWCnJ6x1oX+wD0A3EyjidGXG/kCu8raBuZ7UzwAaWG0fP1jswt
dV/GVE7YCjCagyRrO6fp2rXbQqq4qyZir9nSvHU+h2n9a4mHUD3RBxkQpVVCs9+N
guHQjl4oIBl9vpsB8KyluXdwdrzykk053ryWI7WmwjJdybnUlEShb/w7v359n+Me
DJc9Bd20eDBAB9xJFV8u8gj5Wu13LeacNRHpOz8KcbIfpb2di5MbFjwhaTaXCn/X
4UvR8Sbf+sTR9P1hM1Hrfw0XK570ujC4obqoh93+we4RGkH2s7RZkmzSQmlyWPpb
hqa+hVnHDlOFdinVYfztchbh/lN9xVXnP2zhJFAyceFSgFF9TJUVeUvA8Uqo6w4P
+J7kK0fb9kBfLP7GYVcuknX7lqdGXS0/yjC26ElnqTIg7OfX3lf2OSdx8Xxan7I8
Ps2l3MfClTK2WgNAo6BZiCj32mrj4bi2HWBBlv/CXDAcQ9e1wxgOLJSxYTFAoVYp
8vTZSKweUPSMbr+zbqNCPZZeF4ib93xBQqFBs9o0+bQcT/xMO+5hJTE5GKE07ZG8
5e3QinpBoedoqyz8H8LxwooROqgr0QR6PiVnXGwOekTjUYWx4NXJNw9OQuBT30b+
YpdeNcPSOSqjiybklyoxl46E1fyVMkeL09E9PVTtcQQji5Ts894k4VIDmkIzs+Al
HvRHdYufCUV19kACjShQiGhDz0f9q0OHWf1AuL9+v8wIfnYO5Qy05xAbWNnTVJ6Z
PlP3tj4Dl3hAzU8h+RFgV9U85o24GH8sJDXNpT26LdS14S5IqB5C7VAPFzc+rV3a
c3Mjpyi/QI/w5WV2ngvgQvZR3JbKCCjtyc17n7nrkKNMQb1Copv+aPtUyWEH3AHd
VGsc2EvysmoOa2YYA+0L+cPmAJvxHzyS+8UvpPd23GB0d4e/VKYsH+Ovdz1LfFXd
XhBhINK9tqrKCvVD0MV7wRq5P2dDVePjQ6qdCE/uybajyzd2j6w/Q85mvUbmgTJy
meLfArOISIxkwG/U21ylrZVvQBxJpkHaQVCHho8XmKrBTveZnggNTrrOc2xxkb0p
g2MPPnjOKMEg5xr3XSGpyngo0YSvyv0CENh/XPIpCyOVnTvoow5xrTxn3bpPYyD1
sN05hqzCwQMpcJ0I4fsOpMMeQk7pZ/KW+V/MekSJSrp69ruu2Ri6OoGKKtRnMiRC
JOFzalI/VvhkknO/auDsACec/fjVvOLS2CG1i3E/cJrsxVEgTUgW2x10K89h/Uwz
NLG6vcJBMLT8B+7Ncry0LSZ58PMy7JQGHKUutwSh7qJOhPMlh9RZRd5sJT+tTpRi
s8+136YQrW6yZK60+W9eCGACAC+SQbT5hPCbzT+JxCDtViAFOQO5EhsB33m67gsO
W1DB7ggYjo78Y6XrcW/5CFC/B4ow4oZPY2uVqZLack1Wbg6uw5MDKE4HjML5opoh
Q+Uj+GwLKAsneme9chsV5OjMrFVuB6w8A8oJdI8z9KR5qJqbjZcTztAzqkhyZKuA
LK++lbiqk/EuU4RY/NdQiJ86BzGhkiii2PjKNmqnO6GiTKM8dQyYWccwiL8pjAml
wFnXtxHpONWGDZlUBCcVJX/QewJo0GZObhYqR9K9HvdbwX+JZ5RdqrCOrrrmqXFL
dkVkZOkUgCyudpgWyaLgaQ/S0JlWmfk02boLXmde+DlyPk5Ry8Rvvd8ZKuBm6FFh
LK5vz6kgYldvR2dGl8OCp10g5P8qCZfx+0xJpf/TgEsK8ARYT8rj5Bd6Bt8R2mqT
+QwrI5VQMFCrIqt788lqf/cj+pBKyn8A5KGLyalKrMXUxYWQye8yoxjMRTv4UYaP
NPMbfqbx5voS7fv7OCucd6K7GoYFm99ukEr9eyVVZoKG84PPDpNCz5E9zpBFWEIG
FfmYfxviHX/PA9S5qg9TdYTT0WcLCvIN6HAYb7ROdW1pKe4tdldHdwf0q4A9Fw43
iGOvd7l9iZe4pMXJTF/KFVQM8I6BGYIIZYGkXh0vMm7UN9Lb7SBK73JLcZ+4rdeE
uy6DA0DgV39ccWkQwlupr3dVMghB1vu33mj/SQW0k3qbUV6iNCvV5x8/Bg8g8SBp
cyiAM+ETLGANrq8XIYYvVQ==
//pragma protect end_data_block
//pragma protect digest_block
qkrLt5d8YTujJTTaH5U4OjEjgXc=
//pragma protect end_digest_block
//pragma protect end_protected
